module SG90_LUT (
    input       wire                    i_reset,
    input       wire        [11 : 0]    i_duty,
    output      wire        [11 : 0]    o_duty
);

    parameter                           SERVO_NEUTRAL       =   12'd308;
    reg                     [11 : 0]    r_duty_deg_hex;
    always @(*) begin
        if (i_reset) begin
            r_duty_deg_hex = 0;
        end
        else begin
            if (i_duty >  SERVO_NEUTRAL) begin
                case ((i_duty - SERVO_NEUTRAL))
                    1   :   r_duty_deg_hex = 0;
                    2   :   r_duty_deg_hex = 1;
                    3   :   r_duty_deg_hex = 1;
                    4   :   r_duty_deg_hex = 2;
                    5   :   r_duty_deg_hex = 2;
                    6   :   r_duty_deg_hex = 3;
                    7   :   r_duty_deg_hex = 3;
                    8   :   r_duty_deg_hex = 3;
                    9   :   r_duty_deg_hex = 4;
                    10  :   r_duty_deg_hex = 4;
                    11  :   r_duty_deg_hex = 5;
                    12  :   r_duty_deg_hex = 5;
                    13  :   r_duty_deg_hex = 6;
                    14  :   r_duty_deg_hex = 6;
                    15  :   r_duty_deg_hex = 7;
                    16  :   r_duty_deg_hex = 7;
                    17  :   r_duty_deg_hex = 7;
                    18  :   r_duty_deg_hex = 8;
                    19  :   r_duty_deg_hex = 8;
                    20  :   r_duty_deg_hex = 9;
                    21  :   r_duty_deg_hex = 9;
                    22  :   r_duty_deg_hex = 10;
                    23  :   r_duty_deg_hex = 10;
                    24  :   r_duty_deg_hex = 10;
                    25  :   r_duty_deg_hex = 11;
                    26  :   r_duty_deg_hex = 11;
                    27  :   r_duty_deg_hex = 12;
                    28  :   r_duty_deg_hex = 12;
                    29  :   r_duty_deg_hex = 13;
                    30  :   r_duty_deg_hex = 13;
                    31  :   r_duty_deg_hex = 13;
                    32  :   r_duty_deg_hex = 14;
                    33  :   r_duty_deg_hex = 14;
                    34  :   r_duty_deg_hex = 15;
                    35  :   r_duty_deg_hex = 15;
                    36  :   r_duty_deg_hex = 16;
                    37  :   r_duty_deg_hex = 16;
                    38  :   r_duty_deg_hex = 17;
                    39  :   r_duty_deg_hex = 17;
                    40  :   r_duty_deg_hex = 17;
                    41  :   r_duty_deg_hex = 18;
                    42  :   r_duty_deg_hex = 18;
                    43  :   r_duty_deg_hex = 19;
                    44  :   r_duty_deg_hex = 19;
                    45  :   r_duty_deg_hex = 20;
                    46  :   r_duty_deg_hex = 20;
                    47  :   r_duty_deg_hex = 20;
                    48  :   r_duty_deg_hex = 21;
                    49  :   r_duty_deg_hex = 21;
                    50  :   r_duty_deg_hex = 22;
                    51  :   r_duty_deg_hex = 22;
                    52  :   r_duty_deg_hex = 23;
                    53  :   r_duty_deg_hex = 23;
                    54  :   r_duty_deg_hex = 23;
                    55  :   r_duty_deg_hex = 24;
                    56  :   r_duty_deg_hex = 24;
                    57  :   r_duty_deg_hex = 25;
                    58  :   r_duty_deg_hex = 25;
                    59  :   r_duty_deg_hex = 26;
                    60  :   r_duty_deg_hex = 26;
                    61  :   r_duty_deg_hex = 27;
                    62  :   r_duty_deg_hex = 27;
                    63  :   r_duty_deg_hex = 27;
                    64  :   r_duty_deg_hex = 28;
                    65  :   r_duty_deg_hex = 28;
                    66  :   r_duty_deg_hex = 29;
                    67  :   r_duty_deg_hex = 29;
                    68  :   r_duty_deg_hex = 30;
                    69  :   r_duty_deg_hex = 30;
                    70  :   r_duty_deg_hex = 30;
                    71  :   r_duty_deg_hex = 31;
                    72  :   r_duty_deg_hex = 31;
                    73  :   r_duty_deg_hex = 32;
                    74  :   r_duty_deg_hex = 32;
                    75  :   r_duty_deg_hex = 33;
                    76  :   r_duty_deg_hex = 33;
                    77  :   r_duty_deg_hex = 33;
                    78  :   r_duty_deg_hex = 34;
                    79  :   r_duty_deg_hex = 34;
                    80  :   r_duty_deg_hex = 35;
                    81  :   r_duty_deg_hex = 35;
                    82  :   r_duty_deg_hex = 36;
                    83  :   r_duty_deg_hex = 36;
                    84  :   r_duty_deg_hex = 37;
                    85  :   r_duty_deg_hex = 37;
                    86  :   r_duty_deg_hex = 37;
                    87  :   r_duty_deg_hex = 38;
                    88  :   r_duty_deg_hex = 38;
                    89  :   r_duty_deg_hex = 39;
                    90  :   r_duty_deg_hex = 39;
                    91  :   r_duty_deg_hex = 40;
                    92  :   r_duty_deg_hex = 40;
                    93  :   r_duty_deg_hex = 40;
                    94  :   r_duty_deg_hex = 41;
                    95  :   r_duty_deg_hex = 41;
                    96  :   r_duty_deg_hex = 42;
                    97  :   r_duty_deg_hex = 42;
                    98  :   r_duty_deg_hex = 43;
                    99  :   r_duty_deg_hex = 43;
                    100 :   r_duty_deg_hex = 43;
                    101 :   r_duty_deg_hex = 44;
                    102 :   r_duty_deg_hex = 44;
                    103 :   r_duty_deg_hex = 45;
                    104 :   r_duty_deg_hex = 45;
                    105 :   r_duty_deg_hex = 46;
                    106 :   r_duty_deg_hex = 46;
                    107 :   r_duty_deg_hex = 47;
                    108 :   r_duty_deg_hex = 47;
                    109 :   r_duty_deg_hex = 47;
                    110 :   r_duty_deg_hex = 48;
                    111 :   r_duty_deg_hex = 48;
                    112 :   r_duty_deg_hex = 49;
                    113 :   r_duty_deg_hex = 49;
                    114 :   r_duty_deg_hex = 50;
                    115 :   r_duty_deg_hex = 50;
                    116 :   r_duty_deg_hex = 50;
                    117 :   r_duty_deg_hex = 51;
                    118 :   r_duty_deg_hex = 51;
                    119 :   r_duty_deg_hex = 52;
                    120 :   r_duty_deg_hex = 52;
                    121 :   r_duty_deg_hex = 53;
                    122 :   r_duty_deg_hex = 53;
                    123 :   r_duty_deg_hex = 53;
                    124 :   r_duty_deg_hex = 54;
                    125 :   r_duty_deg_hex = 54;
                    126 :   r_duty_deg_hex = 55;
                    127 :   r_duty_deg_hex = 55;
                    128 :   r_duty_deg_hex = 56;
                    129 :   r_duty_deg_hex = 56;
                    130 :   r_duty_deg_hex = 57;
                    131 :   r_duty_deg_hex = 57;
                    132 :   r_duty_deg_hex = 57;
                    133 :   r_duty_deg_hex = 58;
                    134 :   r_duty_deg_hex = 58;
                    135 :   r_duty_deg_hex = 59;
                    136 :   r_duty_deg_hex = 59;
                    137 :   r_duty_deg_hex = 60;
                    138 :   r_duty_deg_hex = 60;
                    139 :   r_duty_deg_hex = 60;
                    140 :   r_duty_deg_hex = 61;
                    141 :   r_duty_deg_hex = 61;
                    142 :   r_duty_deg_hex = 62;
                    143 :   r_duty_deg_hex = 62;
                    144 :   r_duty_deg_hex = 63;
                    145 :   r_duty_deg_hex = 63;
                    146 :   r_duty_deg_hex = 63;
                    147 :   r_duty_deg_hex = 64;
                    148 :   r_duty_deg_hex = 64;
                    149 :   r_duty_deg_hex = 65;
                    150 :   r_duty_deg_hex = 65;
                    151 :   r_duty_deg_hex = 66;
                    152 :   r_duty_deg_hex = 66;
                    153 :   r_duty_deg_hex = 67;
                    154 :   r_duty_deg_hex = 67;
                    155 :   r_duty_deg_hex = 67;
                    156 :   r_duty_deg_hex = 68;
                    157 :   r_duty_deg_hex = 68;
                    158 :   r_duty_deg_hex = 69;
                    159 :   r_duty_deg_hex = 69;
                    160 :   r_duty_deg_hex = 70;
                    161 :   r_duty_deg_hex = 70;
                    162 :   r_duty_deg_hex = 70;
                    163 :   r_duty_deg_hex = 71;
                    164 :   r_duty_deg_hex = 71;
                    165 :   r_duty_deg_hex = 72;
                    166 :   r_duty_deg_hex = 72;
                    167 :   r_duty_deg_hex = 73;
                    168 :   r_duty_deg_hex = 73;
                    169 :   r_duty_deg_hex = 73;
                    170 :   r_duty_deg_hex = 74;
                    171 :   r_duty_deg_hex = 74;
                    172 :   r_duty_deg_hex = 75;
                    173 :   r_duty_deg_hex = 75;
                    174 :   r_duty_deg_hex = 76;
                    175 :   r_duty_deg_hex = 76;
                    176 :   r_duty_deg_hex = 77;
                    177 :   r_duty_deg_hex = 77;
                    178 :   r_duty_deg_hex = 77;
                    179 :   r_duty_deg_hex = 78;
                    180 :   r_duty_deg_hex = 78;
                    181 :   r_duty_deg_hex = 79;
                    182 :   r_duty_deg_hex = 79;
                    183 :   r_duty_deg_hex = 80;
                    184 :   r_duty_deg_hex = 80;
                    185 :   r_duty_deg_hex = 80;
                    186 :   r_duty_deg_hex = 81;
                    187 :   r_duty_deg_hex = 81;
                    188 :   r_duty_deg_hex = 82;
                    189 :   r_duty_deg_hex = 82;
                    190 :   r_duty_deg_hex = 83;
                    191 :   r_duty_deg_hex = 83;
                    192 :   r_duty_deg_hex = 83;
                    193 :   r_duty_deg_hex = 84;
                    194 :   r_duty_deg_hex = 84;
                    195 :   r_duty_deg_hex = 85;
                    196 :   r_duty_deg_hex = 85;
                    197 :   r_duty_deg_hex = 86;
                    198 :   r_duty_deg_hex = 86;
                    199 :   r_duty_deg_hex = 87;
                    200 :   r_duty_deg_hex = 87;
                    201 :   r_duty_deg_hex = 87;
                    202 :   r_duty_deg_hex = 88;
                    203 :   r_duty_deg_hex = 88;
                    204 :   r_duty_deg_hex = 89;
                    205 :   r_duty_deg_hex = 89;
                    206 :   r_duty_deg_hex = 90;
                    207 :   r_duty_deg_hex = 90;
                    default:r_duty_deg_hex = 0;
                endcase
            end
            else if (i_duty <  SERVO_NEUTRAL) begin
                case ((SERVO_NEUTRAL - i_duty))
                    1   :   r_duty_deg_hex = 0;
                    2   :   r_duty_deg_hex = 1;
                    3   :   r_duty_deg_hex = 1;
                    4   :   r_duty_deg_hex = 2;
                    5   :   r_duty_deg_hex = 2;
                    6   :   r_duty_deg_hex = 3;
                    7   :   r_duty_deg_hex = 3;
                    8   :   r_duty_deg_hex = 3;
                    9   :   r_duty_deg_hex = 4;
                    10  :   r_duty_deg_hex = 4;
                    11  :   r_duty_deg_hex = 5;
                    12  :   r_duty_deg_hex = 5;
                    13  :   r_duty_deg_hex = 6;
                    14  :   r_duty_deg_hex = 6;
                    15  :   r_duty_deg_hex = 7;
                    16  :   r_duty_deg_hex = 7;
                    17  :   r_duty_deg_hex = 7;
                    18  :   r_duty_deg_hex = 8;
                    19  :   r_duty_deg_hex = 8;
                    20  :   r_duty_deg_hex = 9;
                    21  :   r_duty_deg_hex = 9;
                    22  :   r_duty_deg_hex = 10;
                    23  :   r_duty_deg_hex = 10;
                    24  :   r_duty_deg_hex = 10;
                    25  :   r_duty_deg_hex = 11;
                    26  :   r_duty_deg_hex = 11;
                    27  :   r_duty_deg_hex = 12;
                    28  :   r_duty_deg_hex = 12;
                    29  :   r_duty_deg_hex = 13;
                    30  :   r_duty_deg_hex = 13;
                    31  :   r_duty_deg_hex = 13;
                    32  :   r_duty_deg_hex = 14;
                    33  :   r_duty_deg_hex = 14;
                    34  :   r_duty_deg_hex = 15;
                    35  :   r_duty_deg_hex = 15;
                    36  :   r_duty_deg_hex = 16;
                    37  :   r_duty_deg_hex = 16;
                    38  :   r_duty_deg_hex = 17;
                    39  :   r_duty_deg_hex = 17;
                    40  :   r_duty_deg_hex = 17;
                    41  :   r_duty_deg_hex = 18;
                    42  :   r_duty_deg_hex = 18;
                    43  :   r_duty_deg_hex = 19;
                    44  :   r_duty_deg_hex = 19;
                    45  :   r_duty_deg_hex = 20;
                    46  :   r_duty_deg_hex = 20;
                    47  :   r_duty_deg_hex = 20;
                    48  :   r_duty_deg_hex = 21;
                    49  :   r_duty_deg_hex = 21;
                    50  :   r_duty_deg_hex = 22;
                    51  :   r_duty_deg_hex = 22;
                    52  :   r_duty_deg_hex = 23;
                    53  :   r_duty_deg_hex = 23;
                    54  :   r_duty_deg_hex = 23;
                    55  :   r_duty_deg_hex = 24;
                    56  :   r_duty_deg_hex = 24;
                    57  :   r_duty_deg_hex = 25;
                    58  :   r_duty_deg_hex = 25;
                    59  :   r_duty_deg_hex = 26;
                    60  :   r_duty_deg_hex = 26;
                    61  :   r_duty_deg_hex = 27;
                    62  :   r_duty_deg_hex = 27;
                    63  :   r_duty_deg_hex = 27;
                    64  :   r_duty_deg_hex = 28;
                    65  :   r_duty_deg_hex = 28;
                    66  :   r_duty_deg_hex = 29;
                    67  :   r_duty_deg_hex = 29;
                    68  :   r_duty_deg_hex = 30;
                    69  :   r_duty_deg_hex = 30;
                    70  :   r_duty_deg_hex = 30;
                    71  :   r_duty_deg_hex = 31;
                    72  :   r_duty_deg_hex = 31;
                    73  :   r_duty_deg_hex = 32;
                    74  :   r_duty_deg_hex = 32;
                    75  :   r_duty_deg_hex = 33;
                    76  :   r_duty_deg_hex = 33;
                    77  :   r_duty_deg_hex = 33;
                    78  :   r_duty_deg_hex = 34;
                    79  :   r_duty_deg_hex = 34;
                    80  :   r_duty_deg_hex = 35;
                    81  :   r_duty_deg_hex = 35;
                    82  :   r_duty_deg_hex = 36;
                    83  :   r_duty_deg_hex = 36;
                    84  :   r_duty_deg_hex = 37;
                    85  :   r_duty_deg_hex = 37;
                    86  :   r_duty_deg_hex = 37;
                    87  :   r_duty_deg_hex = 38;
                    88  :   r_duty_deg_hex = 38;
                    89  :   r_duty_deg_hex = 39;
                    90  :   r_duty_deg_hex = 39;
                    91  :   r_duty_deg_hex = 40;
                    92  :   r_duty_deg_hex = 40;
                    93  :   r_duty_deg_hex = 40;
                    94  :   r_duty_deg_hex = 41;
                    95  :   r_duty_deg_hex = 41;
                    96  :   r_duty_deg_hex = 42;
                    97  :   r_duty_deg_hex = 42;
                    98  :   r_duty_deg_hex = 43;
                    99  :   r_duty_deg_hex = 43;
                    100 :   r_duty_deg_hex = 43;
                    101 :   r_duty_deg_hex = 44;
                    102 :   r_duty_deg_hex = 44;
                    103 :   r_duty_deg_hex = 45;
                    104 :   r_duty_deg_hex = 45;
                    105 :   r_duty_deg_hex = 46;
                    106 :   r_duty_deg_hex = 46;
                    107 :   r_duty_deg_hex = 47;
                    108 :   r_duty_deg_hex = 47;
                    109 :   r_duty_deg_hex = 47;
                    110 :   r_duty_deg_hex = 48;
                    111 :   r_duty_deg_hex = 48;
                    112 :   r_duty_deg_hex = 49;
                    113 :   r_duty_deg_hex = 49;
                    114 :   r_duty_deg_hex = 50;
                    115 :   r_duty_deg_hex = 50;
                    116 :   r_duty_deg_hex = 50;
                    117 :   r_duty_deg_hex = 51;
                    118 :   r_duty_deg_hex = 51;
                    119 :   r_duty_deg_hex = 52;
                    120 :   r_duty_deg_hex = 52;
                    121 :   r_duty_deg_hex = 53;
                    122 :   r_duty_deg_hex = 53;
                    123 :   r_duty_deg_hex = 53;
                    124 :   r_duty_deg_hex = 54;
                    125 :   r_duty_deg_hex = 54;
                    126 :   r_duty_deg_hex = 55;
                    127 :   r_duty_deg_hex = 55;
                    128 :   r_duty_deg_hex = 56;
                    129 :   r_duty_deg_hex = 56;
                    130 :   r_duty_deg_hex = 57;
                    131 :   r_duty_deg_hex = 57;
                    132 :   r_duty_deg_hex = 57;
                    133 :   r_duty_deg_hex = 58;
                    134 :   r_duty_deg_hex = 58;
                    135 :   r_duty_deg_hex = 59;
                    136 :   r_duty_deg_hex = 59;
                    137 :   r_duty_deg_hex = 60;
                    138 :   r_duty_deg_hex = 60;
                    139 :   r_duty_deg_hex = 60;
                    140 :   r_duty_deg_hex = 61;
                    141 :   r_duty_deg_hex = 61;
                    142 :   r_duty_deg_hex = 62;
                    143 :   r_duty_deg_hex = 62;
                    144 :   r_duty_deg_hex = 63;
                    145 :   r_duty_deg_hex = 63;
                    146 :   r_duty_deg_hex = 63;
                    147 :   r_duty_deg_hex = 64;
                    148 :   r_duty_deg_hex = 64;
                    149 :   r_duty_deg_hex = 65;
                    150 :   r_duty_deg_hex = 65;
                    151 :   r_duty_deg_hex = 66;
                    152 :   r_duty_deg_hex = 66;
                    153 :   r_duty_deg_hex = 67;
                    154 :   r_duty_deg_hex = 67;
                    155 :   r_duty_deg_hex = 67;
                    156 :   r_duty_deg_hex = 68;
                    157 :   r_duty_deg_hex = 68;
                    158 :   r_duty_deg_hex = 69;
                    159 :   r_duty_deg_hex = 69;
                    160 :   r_duty_deg_hex = 70;
                    161 :   r_duty_deg_hex = 70;
                    162 :   r_duty_deg_hex = 70;
                    163 :   r_duty_deg_hex = 71;
                    164 :   r_duty_deg_hex = 71;
                    165 :   r_duty_deg_hex = 72;
                    166 :   r_duty_deg_hex = 72;
                    167 :   r_duty_deg_hex = 73;
                    168 :   r_duty_deg_hex = 73;
                    169 :   r_duty_deg_hex = 73;
                    170 :   r_duty_deg_hex = 74;
                    171 :   r_duty_deg_hex = 74;
                    172 :   r_duty_deg_hex = 75;
                    173 :   r_duty_deg_hex = 75;
                    174 :   r_duty_deg_hex = 76;
                    175 :   r_duty_deg_hex = 76;
                    176 :   r_duty_deg_hex = 77;
                    177 :   r_duty_deg_hex = 77;
                    178 :   r_duty_deg_hex = 77;
                    179 :   r_duty_deg_hex = 78;
                    180 :   r_duty_deg_hex = 78;
                    181 :   r_duty_deg_hex = 79;
                    182 :   r_duty_deg_hex = 79;
                    183 :   r_duty_deg_hex = 80;
                    184 :   r_duty_deg_hex = 80;
                    185 :   r_duty_deg_hex = 80;
                    186 :   r_duty_deg_hex = 81;
                    187 :   r_duty_deg_hex = 81;
                    188 :   r_duty_deg_hex = 82;
                    189 :   r_duty_deg_hex = 82;
                    190 :   r_duty_deg_hex = 83;
                    191 :   r_duty_deg_hex = 83;
                    192 :   r_duty_deg_hex = 83;
                    193 :   r_duty_deg_hex = 84;
                    194 :   r_duty_deg_hex = 84;
                    195 :   r_duty_deg_hex = 85;
                    196 :   r_duty_deg_hex = 85;
                    197 :   r_duty_deg_hex = 86;
                    198 :   r_duty_deg_hex = 86;
                    199 :   r_duty_deg_hex = 87;
                    200 :   r_duty_deg_hex = 87;
                    201 :   r_duty_deg_hex = 87;
                    202 :   r_duty_deg_hex = 88;
                    203 :   r_duty_deg_hex = 88;
                    204 :   r_duty_deg_hex = 89;
                    205 :   r_duty_deg_hex = 89;
                    206 :   r_duty_deg_hex = 90;
                    207 :   r_duty_deg_hex = 90;
                    default:r_duty_deg_hex = 0;
                endcase
            end
            else begin
                r_duty_deg_hex = 0;
            end
        end
    end

    assign o_duty = r_duty_deg_hex;
    
endmodule
//////////////////////////////////////////////////////////////////////////////////
module Q8_8_Mapper (
    input       wire        signed      [7 : 0]         i_binVal,
    output      wire        signed      [15 : 0]        o_qVal
);

    assign o_qVal = i_binVal << 8;

endmodule
//////////////////////////////////////////////////////////////////////////////////
module BIN_Mapper #(
    parameter                           INTEGER_WIDTH   =   16
)(
    input       wire        signed      [2*INTEGER_WIDTH - 1 : 0]        i_qVal,
    output      wire        signed      [INTEGER_WIDTH - 1   : 0]        o_binVal
);

    assign o_binVal = i_qVal[2*INTEGER_WIDTH - 1 -: INTEGER_WIDTH];
    
endmodule

//////////////////////////////////////////////////////////////////////////////////
module sin_LUT (
    input       wire                                    i_reset,
    input       wire        signed      [15 : 0]        i_radVal_q8_8,
    output      wire        signed      [15 : 0]        o_sinVal_q8_8
);
                reg         signed      [15 : 0]        r_sinVal;

    always @(*) begin
        if (i_reset) begin
            r_sinVal = 0;
        end
        else begin
            case (i_radVal_q8_8)
                0   :   r_sinVal = 0;
                1   :   r_sinVal = 1;
                2   :   r_sinVal = 2;
                3   :   r_sinVal = 3;
                4   :   r_sinVal = 4;
                5   :   r_sinVal = 5;
                6   :   r_sinVal = 6;
                7   :   r_sinVal = 7;
                8   :   r_sinVal = 8;
                9   :   r_sinVal = 9;
                10  :   r_sinVal = 10;
                11  :   r_sinVal = 11;
                12  :   r_sinVal = 12;
                13  :   r_sinVal = 13;
                14  :   r_sinVal = 14;
                15  :   r_sinVal = 15;
                16  :   r_sinVal = 16;
                17  :   r_sinVal = 17;
                18  :   r_sinVal = 18;
                19  :   r_sinVal = 19;
                20  :   r_sinVal = 20;
                21  :   r_sinVal = 21;
                22  :   r_sinVal = 22;
                23  :   r_sinVal = 23;
                24  :   r_sinVal = 24;
                25  :   r_sinVal = 25;
                26  :   r_sinVal = 26;
                27  :   r_sinVal = 27;
                28  :   r_sinVal = 28;
                29  :   r_sinVal = 29;
                30  :   r_sinVal = 30;
                31  :   r_sinVal = 31;
                32  :   r_sinVal = 32;
                33  :   r_sinVal = 33;
                34  :   r_sinVal = 34;
                35  :   r_sinVal = 35;
                36  :   r_sinVal = 36;
                37  :   r_sinVal = 37;
                38  :   r_sinVal = 38;
                39  :   r_sinVal = 39;
                40  :   r_sinVal = 40;
                41  :   r_sinVal = 41;
                42  :   r_sinVal = 42;
                43  :   r_sinVal = 43;
                44  :   r_sinVal = 44;
                45  :   r_sinVal = 44;
                46  :   r_sinVal = 46;
                47  :   r_sinVal = 47;
                48  :   r_sinVal = 48;
                49  :   r_sinVal = 49;
                50  :   r_sinVal = 50;
                51  :   r_sinVal = 51;
                52  :   r_sinVal = 52;
                53  :   r_sinVal = 53;
                54  :   r_sinVal = 53;
                55  :   r_sinVal = 55;
                56  :   r_sinVal = 56;
                57  :   r_sinVal = 57;
                58  :   r_sinVal = 58;
                59  :   r_sinVal = 59;
                60  :   r_sinVal = 60;
                61  :   r_sinVal = 61;
                62  :   r_sinVal = 62;
                63  :   r_sinVal = 62;
                63  :   r_sinVal = 62;
                64  :   r_sinVal = 64;
                65  :   r_sinVal = 65;
                66  :   r_sinVal = 66;
                67  :   r_sinVal = 66;
                68  :   r_sinVal = 68;
                69  :   r_sinVal = 69;
                70  :   r_sinVal = 70;
                71  :   r_sinVal = 71;
                72  :   r_sinVal = 72;
                73  :   r_sinVal = 73;
                74  :   r_sinVal = 74;
                75  :   r_sinVal = 75;
                76  :   r_sinVal = 75;
                77  :   r_sinVal = 77;
                78  :   r_sinVal = 78;
                79  :   r_sinVal = 79;
                80  :   r_sinVal = 79;
                81  :   r_sinVal = 80;
                82  :   r_sinVal = 81;
                83  :   r_sinVal = 82;
                84  :   r_sinVal = 83;
                85  :   r_sinVal = 83;
                86  :   r_sinVal = 86;
                87  :   r_sinVal = 87;
                88  :   r_sinVal = 88;
                89  :   r_sinVal = 88;
                90  :   r_sinVal = 90;
                91  :   r_sinVal = 90;
                92  :   r_sinVal = 91;
                93  :   r_sinVal = 91;
                94  :   r_sinVal = 92;
                95  :   r_sinVal = 93;
                96  :   r_sinVal = 94;
                97  :   r_sinVal = 95;
                98  :   r_sinVal = 96;
                99  :   r_sinVal = 97;
                100 :   r_sinVal = 98;
                101 :   r_sinVal = 99;
                102 :   r_sinVal = 100;
                103 :   r_sinVal = 100;
                104 :   r_sinVal = 101;
                105 :   r_sinVal = 102;
                106 :   r_sinVal = 103;
                107 :   r_sinVal = 104;
                108 :   r_sinVal = 104;
                109 :   r_sinVal = 105;
                110 :   r_sinVal = 106;
                111 :   r_sinVal = 107;
                112 :   r_sinVal = 108;
                113 :   r_sinVal = 109;
                114 :   r_sinVal = 110;
                115 :   r_sinVal = 111;
                116 :   r_sinVal = 111;
                117 :   r_sinVal = 112;
                118 :   r_sinVal = 113;
                119 :   r_sinVal = 114;
                120 :   r_sinVal = 115;
                121 :   r_sinVal = 116;
                125 :   r_sinVal = 120;
                126 :   r_sinVal = 120;
                127 :   r_sinVal = 121;
                128 :   r_sinVal = 122;
                129 :   r_sinVal = 123;
                130 :   r_sinVal = 124;
                131 :   r_sinVal = 125;
                132 :   r_sinVal = 126;
                133 :   r_sinVal = 127;
                134 :   r_sinVal = 128;
                135 :   r_sinVal = 128;
                136 :   r_sinVal = 129;
                137 :   r_sinVal = 130;
                138 :   r_sinVal = 131;
                139 :   r_sinVal = 132;
                140 :   r_sinVal = 133;
                141 :   r_sinVal = 134;
                142 :   r_sinVal = 135;
                143 :   r_sinVal = 136;
                144 :   r_sinVal = 136;
                145 :   r_sinVal = 137;
                146 :   r_sinVal = 138;
                147 :   r_sinVal = 139;
                148 :   r_sinVal = 139;
                149 :   r_sinVal = 140;
                150 :   r_sinVal = 141;
                151 :   r_sinVal = 142;
                152 :   r_sinVal = 143;
                153 :   r_sinVal = 144;
                154 :   r_sinVal = 145;
                155 :   r_sinVal = 146;
                156 :   r_sinVal = 147;
                157 :   r_sinVal = 147;
                158 :   r_sinVal = 147;
                159 :   r_sinVal = 148;
                160 :   r_sinVal = 149;
                161 :   r_sinVal = 150;
                162 :   r_sinVal = 151;
                163 :   r_sinVal = 152;
                164 :   r_sinVal = 153;
                165 :   r_sinVal = 154;
                166 :   r_sinVal = 154;
                167 :   r_sinVal = 155;
                168 :   r_sinVal = 156;
                169 :   r_sinVal = 157;
                170 :   r_sinVal = 158;
                171 :   r_sinVal = 158;
                172 :   r_sinVal = 159;
                173 :   r_sinVal = 160;
                174 :   r_sinVal = 161;
                175 :   r_sinVal = 161;
                176 :   r_sinVal = 162;
                177 :   r_sinVal = 163;
                178 :   r_sinVal = 164;
                179 :   r_sinVal = 164;
                180 :   r_sinVal = 165;
                181 :   r_sinVal = 166;
                182 :   r_sinVal = 167;
                183 :   r_sinVal = 167;
                184 :   r_sinVal = 168;
                185 :   r_sinVal = 168;
                186 :   r_sinVal = 169;
                187 :   r_sinVal = 170;
                188 :   r_sinVal = 171;
                189 :   r_sinVal = 172;
                190 :   r_sinVal = 173;
                191 :   r_sinVal = 174;
                192 :   r_sinVal = 174;
                193 :   r_sinVal = 175;
                194 :   r_sinVal = 175;
                195 :   r_sinVal = 176;
                196 :   r_sinVal = 177;
                197 :   r_sinVal = 178;
                198 :   r_sinVal = 179;
                199 :   r_sinVal = 180;
                200 :   r_sinVal = 180;
                201 :   r_sinVal = 181;
                202 :   r_sinVal = 181;
                203 :   r_sinVal = 182;
                204 :   r_sinVal = 182;
                205 :   r_sinVal = 183;
                206 :   r_sinVal = 184;
                207 :   r_sinVal = 184;
                208 :   r_sinVal = 185;
                209 :   r_sinVal = 186;
                210 :   r_sinVal = 187;
                211 :   r_sinVal = 187;
                212 :   r_sinVal = 188;
                213 :   r_sinVal = 189;
                214 :   r_sinVal = 190;
                215 :   r_sinVal = 191;
                216 :   r_sinVal = 191;
                217 :   r_sinVal = 192;
                218 :   r_sinVal = 192;
                219 :   r_sinVal = 193;
                220 :   r_sinVal = 193;
                221 :   r_sinVal = 194;
                222 :   r_sinVal = 195;
                223 :   r_sinVal = 195;
                224 :   r_sinVal = 196;
                225 :   r_sinVal = 197;
                226 :   r_sinVal = 197;
                227 :   r_sinVal = 198;
                228 :   r_sinVal = 199;
                229 :   r_sinVal = 200;
                230 :   r_sinVal = 201;
                231 :   r_sinVal = 202;
                232 :   r_sinVal = 202;
                233 :   r_sinVal = 203;
                234 :   r_sinVal = 203;
                235 :   r_sinVal = 204;
                236 :   r_sinVal = 204;
                237 :   r_sinVal = 205;
                238 :   r_sinVal = 205;
                239 :   r_sinVal = 206;
                240 :   r_sinVal = 207;
                241 :   r_sinVal = 207;
                242 :   r_sinVal = 208;
                243 :   r_sinVal = 208;
                244 :   r_sinVal = 209;
                245 :   r_sinVal = 210;
                246 :   r_sinVal = 210;
                247 :   r_sinVal = 211;
                248 :   r_sinVal = 211;
                249 :   r_sinVal = 212;
                250 :   r_sinVal = 212;
                251 :   r_sinVal = 213;
                252 :   r_sinVal = 213;
                253 :   r_sinVal = 214;
                254 :   r_sinVal = 215;
                255 :   r_sinVal = 215;
                256 :   r_sinVal = 216;
                257 :   r_sinVal = 216;
                258 :   r_sinVal = 217;
                259 :   r_sinVal = 217;
                260 :   r_sinVal = 217;
                261 :   r_sinVal = 218;
                262 :   r_sinVal = 218;
                263 :   r_sinVal = 219;
                264 :   r_sinVal = 219;
                265 :   r_sinVal = 220;
                266 :   r_sinVal = 220;
                267 :   r_sinVal = 221;
                268 :   r_sinVal = 222;
                269 :   r_sinVal = 222;
                270 :   r_sinVal = 223;
                271 :   r_sinVal = 223;
                272 :   r_sinVal = 224;
                273 :   r_sinVal = 224;
                274 :   r_sinVal = 225;
                275 :   r_sinVal = 225;
                276 :   r_sinVal = 226;
                277 :   r_sinVal = 226;
                278 :   r_sinVal = 227;
                279 :   r_sinVal = 227;
                280 :   r_sinVal = 228;
                281 :   r_sinVal = 228;
                282 :   r_sinVal = 228;
                283 :   r_sinVal = 229;
                284 :   r_sinVal = 229;
                285 :   r_sinVal = 230;
                286 :   r_sinVal = 230;
                287 :   r_sinVal = 231;
                288 :   r_sinVal = 231;
                289 :   r_sinVal = 232;
                290 :   r_sinVal = 232;
                291 :   r_sinVal = 232;
                292 :   r_sinVal = 233;
                293 :   r_sinVal = 233;
                294 :   r_sinVal = 234;
                295 :   r_sinVal = 234;
                296 :   r_sinVal = 235;
                297 :   r_sinVal = 235;
                298 :   r_sinVal = 236;
                299 :   r_sinVal = 236;
                300 :   r_sinVal = 236;
                301 :   r_sinVal = 236;
                302 :   r_sinVal = 236;
                303 :   r_sinVal = 237;
                304 :   r_sinVal = 237;
                305 :   r_sinVal = 238;
                306 :   r_sinVal = 238;
                307 :   r_sinVal = 239;
                308 :   r_sinVal = 239;
                309 :   r_sinVal = 239;
                310 :   r_sinVal = 240;
                311 :   r_sinVal = 240;
                312 :   r_sinVal = 241;
                313 :   r_sinVal = 241;
                314 :   r_sinVal = 241;
                315 :   r_sinVal = 242;
                316 :   r_sinVal = 242;
                317 :   r_sinVal = 242;
                318 :   r_sinVal = 242;
                319 :   r_sinVal = 242;
                320 :   r_sinVal = 242;
                321 :   r_sinVal = 243;
                322 :   r_sinVal = 243;
                323 :   r_sinVal = 244;
                324 :   r_sinVal = 244;
                325 :   r_sinVal = 245;
                326 :   r_sinVal = 245;
                327 :   r_sinVal = 245;
                328 :   r_sinVal = 245;
                329 :   r_sinVal = 246;
                330 :   r_sinVal = 246;
                331 :   r_sinVal = 246;
                332 :   r_sinVal = 246;
                333 :   r_sinVal = 247;
                334 :   r_sinVal = 247;
                335 :   r_sinVal = 247;
                336 :   r_sinVal = 247;
                337 :   r_sinVal = 248;
                338 :   r_sinVal = 248;
                339 :   r_sinVal = 248;
                340 :   r_sinVal = 248;
                341 :   r_sinVal = 248;
                342 :   r_sinVal = 249;
                343 :   r_sinVal = 249;
                344 :   r_sinVal = 249;
                345 :   r_sinVal = 249;
                346 :   r_sinVal = 250;
                347 :   r_sinVal = 250;
                348 :   r_sinVal = 250;
                349 :   r_sinVal = 250;
                350 :   r_sinVal = 251;
                351 :   r_sinVal = 251;
                352 :   r_sinVal = 251;
                353 :   r_sinVal = 251;
                354 :   r_sinVal = 252;
                355 :   r_sinVal = 252;
                356 :   r_sinVal = 252;
                357 :   r_sinVal = 252;
                358 :   r_sinVal = 253;
                359 :   r_sinVal = 253;
                360 :   r_sinVal = 253;
                361 :   r_sinVal = 253;
                362 :   r_sinVal = 253;
                363 :   r_sinVal = 254;
                364 :   r_sinVal = 254;
                365 :   r_sinVal = 254;
                366 :   r_sinVal = 254;
                367 :   r_sinVal = 254;
                368 :   r_sinVal = 254;
                369 :   r_sinVal = 254;
                370 :   r_sinVal = 254;
                371 :   r_sinVal = 255;
                372 :   r_sinVal = 255;
                373 :   r_sinVal = 255;
                374 :   r_sinVal = 255;
                375 :   r_sinVal = 255;
                376 :   r_sinVal = 255;
                377 :   r_sinVal = 255;
                378 :   r_sinVal = 255;
                379 :   r_sinVal = 255;
                380 :   r_sinVal = 255;
                384 :   r_sinVal = 255;
                385 :   r_sinVal = 255;
                386 :   r_sinVal = 256;
                387 :   r_sinVal = 256;
                388 :   r_sinVal = 256;
                389 :   r_sinVal = 256;
                390 :   r_sinVal = 256;
                391 :   r_sinVal = 256;
                392 :   r_sinVal = 256;
                393 :   r_sinVal = 256;
                394 :   r_sinVal = 256;
                395 :   r_sinVal = 256;
                396 :   r_sinVal = 256;
                397 :   r_sinVal = 256;
                398 :   r_sinVal = 256;
                399 :   r_sinVal = 256;
                400 :   r_sinVal = 256;
                401 :   r_sinVal = 256;
                402 :   r_sinVal = 256;
                403 :   r_sinVal = 256;
                404 :   r_sinVal = 256;
                405 :   r_sinVal = 256;
                406 :   r_sinVal = 256;
                407 :   r_sinVal = 256;
                408 :   r_sinVal = 256;
                409 :   r_sinVal = 256;
                410 :   r_sinVal = 256;
                411 :   r_sinVal = 256;
                412 :   r_sinVal = 256;
                413 :   r_sinVal = 256;
                414 :   r_sinVal = 256;
                415 :   r_sinVal = 256;
                416 :   r_sinVal = 256;
                420 :   r_sinVal = 255;
                421 :   r_sinVal = 255;
                422 :   r_sinVal = 255;
                423 :   r_sinVal = 255;
                424 :   r_sinVal = 255;
                425 :   r_sinVal = 255;
                426 :   r_sinVal = 255;
                427 :   r_sinVal = 255;
                428 :   r_sinVal = 255;
                429 :   r_sinVal = 255;
                430 :   r_sinVal = 254;
                431 :   r_sinVal = 254;
                432 :   r_sinVal = 254;
                433 :   r_sinVal = 254;
                434 :   r_sinVal = 254;
                435 :   r_sinVal = 254;
                436 :   r_sinVal = 254;
                437 :   r_sinVal = 254;
                438 :   r_sinVal = 253;
                439 :   r_sinVal = 253;
                440 :   r_sinVal = 253;
                441 :   r_sinVal = 253;
                442 :   r_sinVal = 253;
                443 :   r_sinVal = 252;
                444 :   r_sinVal = 252;
                445 :   r_sinVal = 252;
                446 :   r_sinVal = 252;
                447 :   r_sinVal = 251;
                448 :   r_sinVal = 251;
                449 :   r_sinVal = 251;
                450 :   r_sinVal = 251;
                451 :   r_sinVal = 251;
                452 :   r_sinVal = 251;
                453 :   r_sinVal = 250;
                454 :   r_sinVal = 250;
                455 :   r_sinVal = 250;
                456 :   r_sinVal = 250;
                457 :   r_sinVal = 249;
                458 :   r_sinVal = 249;
                459 :   r_sinVal = 249;
                460 :   r_sinVal = 249;
                461 :   r_sinVal = 249;
                462 :   r_sinVal = 248;
                463 :   r_sinVal = 248;
                464 :   r_sinVal = 248;
                465 :   r_sinVal = 248;
                466 :   r_sinVal = 247;
                467 :   r_sinVal = 247;
                468 :   r_sinVal = 247;
                469 :   r_sinVal = 247;
                470 :   r_sinVal = 247;
                471 :   r_sinVal = 246;
                472 :   r_sinVal = 246;
                473 :   r_sinVal = 246;
                474 :   r_sinVal = 246;
                475 :   r_sinVal = 245;
                476 :   r_sinVal = 245;
                477 :   r_sinVal = 245;
                478 :   r_sinVal = 245;
                479 :   r_sinVal = 244;
                480 :   r_sinVal = 244;
                481 :   r_sinVal = 244;
                482 :   r_sinVal = 244;
                483 :   r_sinVal = 243;
                484 :   r_sinVal = 243;
                485 :   r_sinVal = 243;
                486 :   r_sinVal = 242;
                487 :   r_sinVal = 242;
                488 :   r_sinVal = 242;
                489 :   r_sinVal = 241;
                490 :   r_sinVal = 241;
                491 :   r_sinVal = 241;
                492 :   r_sinVal = 241;
                493 :   r_sinVal = 240;
                494 :   r_sinVal = 240;
                495 :   r_sinVal = 240;
                496 :   r_sinVal = 239;
                497 :   r_sinVal = 239;
                498 :   r_sinVal = 239;
                499 :   r_sinVal = 239;
                500 :   r_sinVal = 238;
                501 :   r_sinVal = 238;
                502 :   r_sinVal = 238;
                503 :   r_sinVal = 237;
                504 :   r_sinVal = 237;
                505 :   r_sinVal = 236;
                506 :   r_sinVal = 236;
                507 :   r_sinVal = 235;
                508 :   r_sinVal = 235;
                509 :   r_sinVal = 234;
                510 :   r_sinVal = 234;
                511 :   r_sinVal = 234;
                512 :   r_sinVal = 233;
                513 :   r_sinVal = 233;
                514 :   r_sinVal = 232;
                515 :   r_sinVal = 232;
                516 :   r_sinVal = 231;
                517 :   r_sinVal = 231;
                518 :   r_sinVal = 230;
                519 :   r_sinVal = 230;
                520 :   r_sinVal = 229;
                521 :   r_sinVal = 229;
                522 :   r_sinVal = 229;
                523 :   r_sinVal = 228;
                524 :   r_sinVal = 228;
                525 :   r_sinVal = 227;
                526 :   r_sinVal = 227;
                527 :   r_sinVal = 226;
                528 :   r_sinVal = 226;
                529 :   r_sinVal = 226;
                530 :   r_sinVal = 225;
                531 :   r_sinVal = 225;
                532 :   r_sinVal = 224;
                533 :   r_sinVal = 224;
                534 :   r_sinVal = 223;
                535 :   r_sinVal = 223;
                536 :   r_sinVal = 222;
                537 :   r_sinVal = 222;
                538 :   r_sinVal = 221;
                539 :   r_sinVal = 221;
                540 :   r_sinVal = 220;
                541 :   r_sinVal = 220;
                542 :   r_sinVal = 219;
                543 :   r_sinVal = 219;
                544 :   r_sinVal = 218;
                545 :   r_sinVal = 217;
                546 :   r_sinVal = 217;
                547 :   r_sinVal = 217;
                548 :   r_sinVal = 216;
                549 :   r_sinVal = 216;
                550 :   r_sinVal = 215;
                551 :   r_sinVal = 215;
                552 :   r_sinVal = 214;
                553 :   r_sinVal = 213;
                554 :   r_sinVal = 212;
                555 :   r_sinVal = 212;
                556 :   r_sinVal = 212;
                557 :   r_sinVal = 211;
                558 :   r_sinVal = 211;
                559 :   r_sinVal = 210;
                560 :   r_sinVal = 209;
                561 :   r_sinVal = 208;
                562 :   r_sinVal = 207;
                563 :   r_sinVal = 207;
                564 :   r_sinVal = 206;
                565 :   r_sinVal = 205;
                566 :   r_sinVal = 205;
                567 :   r_sinVal = 204;
                568 :   r_sinVal = 204;
                569 :   r_sinVal = 203;
                570 :   r_sinVal = 203;
                571 :   r_sinVal = 202;
                572 :   r_sinVal = 202;
                573 :   r_sinVal = 201;
                574 :   r_sinVal = 201;
                575 :   r_sinVal = 200;
                576 :   r_sinVal = 199;
                577 :   r_sinVal = 199;
                578 :   r_sinVal = 198;
                579 :   r_sinVal = 198;
                580 :   r_sinVal = 197;
                581 :   r_sinVal = 196;
                582 :   r_sinVal = 195;
                583 :   r_sinVal = 194;
                584 :   r_sinVal = 193;
                585 :   r_sinVal = 193;
                586 :   r_sinVal = 192;
                587 :   r_sinVal = 192;
                588 :   r_sinVal = 191;
                589 :   r_sinVal = 191;
                590 :   r_sinVal = 190;
                591 :   r_sinVal = 190;
                592 :   r_sinVal = 189;
                593 :   r_sinVal = 188;
                594 :   r_sinVal = 187;
                595 :   r_sinVal = 187;
                596 :   r_sinVal = 186;
                597 :   r_sinVal = 185;
                598 :   r_sinVal = 185;
                599 :   r_sinVal = 184;
                600 :   r_sinVal = 184;
                601 :   r_sinVal = 183;
                602 :   r_sinVal = 182;
                603 :   r_sinVal = 181;
                604 :   r_sinVal = 181;
                605 :   r_sinVal = 180;
                606 :   r_sinVal = 179;
                607 :   r_sinVal = 178;
                608 :   r_sinVal = 178;
                609 :   r_sinVal = 177;
                610 :   r_sinVal = 176;
                611 :   r_sinVal = 175;
                612 :   r_sinVal = 175;
                613 :   r_sinVal = 174;
                614 :   r_sinVal = 174;
                615 :   r_sinVal = 173;
                616 :   r_sinVal = 172;
                617 :   r_sinVal = 171;
                618 :   r_sinVal = 170;
                619 :   r_sinVal = 169;
                620 :   r_sinVal = 168;
                621 :   r_sinVal = 168;
                622 :   r_sinVal = 167;
                623 :   r_sinVal = 166;
                624 :   r_sinVal = 166;
                625 :   r_sinVal = 165;
                626 :   r_sinVal = 165;
                627 :   r_sinVal = 164;
                628 :   r_sinVal = 163;
                629 :   r_sinVal = 162;
                630 :   r_sinVal = 161;
                631 :   r_sinVal = 161;
                632 :   r_sinVal = 160;
                633 :   r_sinVal = 159;
                634 :   r_sinVal = 158;
                635 :   r_sinVal = 158;
                636 :   r_sinVal = 157;
                637 :   r_sinVal = 156;
                638 :   r_sinVal = 155;
                639 :   r_sinVal = 154;
                640 :   r_sinVal = 153;
                641 :   r_sinVal = 152;
                642 :   r_sinVal = 151;
                643 :   r_sinVal = 150;
                644 :   r_sinVal = 150;
                645 :   r_sinVal = 150;
                646 :   r_sinVal = 149;
                647 :   r_sinVal = 148;
                648 :   r_sinVal = 147;
                649 :   r_sinVal = 146;
                650 :   r_sinVal = 145;
                651 :   r_sinVal = 144;
                652 :   r_sinVal = 143;
                653 :   r_sinVal = 142;
                654 :   r_sinVal = 141;
                655 :   r_sinVal = 140;
                656 :   r_sinVal = 139;
                657 :   r_sinVal = 139;
                658 :   r_sinVal = 138;
                659 :   r_sinVal = 138;
                660 :   r_sinVal = 137;
                661 :   r_sinVal = 136;
                662 :   r_sinVal = 135;
                663 :   r_sinVal = 134;
                664 :   r_sinVal = 133;
                665 :   r_sinVal = 133;
                666 :   r_sinVal = 132;
                667 :   r_sinVal = 131;
                668 :   r_sinVal = 130;
                669 :   r_sinVal = 129;
                670 :   r_sinVal = 128;
                671 :   r_sinVal = 127;
                672 :   r_sinVal = 126;
                673 :   r_sinVal = 125;
                674 :   r_sinVal = 125;
                675 :   r_sinVal = 124;
                676 :   r_sinVal = 123;
                677 :   r_sinVal = 122;
                678 :   r_sinVal = 121;
                679 :   r_sinVal = 120;
                680 :   r_sinVal = 120;
                681 :   r_sinVal = 119;
                682 :   r_sinVal = 118;
                683 :   r_sinVal = 117;
                684 :   r_sinVal = 116;
                685 :   r_sinVal = 115;
                686 :   r_sinVal = 114;
                687 :   r_sinVal = 113;
                688 :   r_sinVal = 112;
                689 :   r_sinVal = 112;
                690 :   r_sinVal = 111;
                691 :   r_sinVal = 110;
                692 :   r_sinVal = 109;
                693 :   r_sinVal = 108;
                694 :   r_sinVal = 107;
                695 :   r_sinVal = 106;
                696 :   r_sinVal = 105;
                697 :   r_sinVal = 104;
                698 :   r_sinVal = 103;
                699 :   r_sinVal = 102;
                700 :   r_sinVal = 101;
                701 :   r_sinVal = 100;
                702 :   r_sinVal = 100;
                703 :   r_sinVal = 99;
                704 :   r_sinVal = 98;
                705 :   r_sinVal = 97;
                706 :   r_sinVal = 96;
                707 :   r_sinVal = 96;
                708 :   r_sinVal = 95;
                709 :   r_sinVal = 94;
                710 :   r_sinVal = 93;
                711 :   r_sinVal = 92;
                712 :   r_sinVal = 91;
                713 :   r_sinVal = 90;
                714 :   r_sinVal = 89;
                715 :   r_sinVal = 88;
                716 :   r_sinVal = 87;
                717 :   r_sinVal = 86;
                718 :   r_sinVal = 85;
                719 :   r_sinVal = 84;
                720 :   r_sinVal = 83;
                721 :   r_sinVal = 82;
                722 :   r_sinVal = 81;
                723 :   r_sinVal = 80;
                724 :   r_sinVal = 79;
                725 :   r_sinVal = 78;
                726 :   r_sinVal = 77;
                727 :   r_sinVal = 76;
                728 :   r_sinVal = 75;
                729 :   r_sinVal = 74;
                730 :   r_sinVal = 73;
                731 :   r_sinVal = 72;
                732 :   r_sinVal = 71;
                733 :   r_sinVal = 70;
                734 :   r_sinVal = 69;
                735 :   r_sinVal = 68;
                736 :   r_sinVal = 67;
                737 :   r_sinVal = 66;
                738 :   r_sinVal = 65;
                739 :   r_sinVal = 64;
                740 :   r_sinVal = 63;
                741 :   r_sinVal = 62;
                742 :   r_sinVal = 61;
                743 :   r_sinVal = 60;
                744 :   r_sinVal = 59;
                745 :   r_sinVal = 59;
                746 :   r_sinVal = 58;
                747 :   r_sinVal = 57;
                748 :   r_sinVal = 56;
                749 :   r_sinVal = 55;
                750 :   r_sinVal = 54;
                751 :   r_sinVal = 53;
                752 :   r_sinVal = 52;
                753 :   r_sinVal = 51;
                754 :   r_sinVal = 50;
                755 :   r_sinVal = 49;
                756 :   r_sinVal = 48;
                757 :   r_sinVal = 47;
                758 :   r_sinVal = 46;
                759 :   r_sinVal = 45;
                760 :   r_sinVal = 44;
                761 :   r_sinVal = 43;
                762 :   r_sinVal = 42;
                763 :   r_sinVal = 41;
                764 :   r_sinVal = 40;
                765 :   r_sinVal = 39;
                766 :   r_sinVal = 38;
                767 :   r_sinVal = 37;
                768 :   r_sinVal = 36;
                769 :   r_sinVal = 35;
                770 :   r_sinVal = 34;
                771 :   r_sinVal = 33;
                772 :   r_sinVal = 32;
                773 :   r_sinVal = 31;
                774 :   r_sinVal = 30;
                775 :   r_sinVal = 29;
                776 :   r_sinVal = 28;
                777 :   r_sinVal = 27;
                778 :   r_sinVal = 26;
                779 :   r_sinVal = 25;
                780 :   r_sinVal = 24;
                781 :   r_sinVal = 23;
                782 :   r_sinVal = 22;
                783 :   r_sinVal = 21;
                784 :   r_sinVal = 20;
                785 :   r_sinVal = 19;
                786 :   r_sinVal = 18;
                787 :   r_sinVal = 17;
                788 :   r_sinVal = 16;
                789 :   r_sinVal = 15;
                790 :   r_sinVal = 14;
                791 :   r_sinVal = 13;
                792 :   r_sinVal = 12;
                793 :   r_sinVal = 11;
                794 :   r_sinVal = 10;
                795 :   r_sinVal = 9;
                796 :   r_sinVal = 8;
                797 :   r_sinVal = 7;
                798 :   r_sinVal = 6;
                799 :   r_sinVal = 5;
                800 :   r_sinVal = 4;
                800 :   r_sinVal = 3;
                800 :   r_sinVal = 2;
                800 :   r_sinVal = 1;
                804 :   r_sinVal = 0;
                default : r_sinVal = r_sinVal;
            endcase
        end
    end

    assign o_sinVal_q8_8 = r_sinVal;

endmodule
//////////////////////////////////////////////////////////////////////////////////
module cos_LUT (
    input       wire                                    i_reset,
    input       wire        signed      [15 : 0]        i_radVal_q8_8,
    output      wire        signed      [15 : 0]        o_cosVal_q8_8
);
                reg         signed      [15 : 0]        r_cosVal;

    always @(*) begin
        if (i_reset) begin
            r_cosVal = 0;
        end
        else begin
            case (i_radVal_q8_8)
                0   :   r_cosVal = 256;
                4   :   r_cosVal = 256;
                9   :   r_cosVal = 256;
                13  :   r_cosVal = 256;
                18  :   r_cosVal = 255;
                22  :   r_cosVal = 255;
                27  :   r_cosVal = 255;
                31  :   r_cosVal = 254;
                36  :   r_cosVal = 254;
                40  :   r_cosVal = 253;
                45  :   r_cosVal = 252;
                49  :   r_cosVal = 251;
                54  :   r_cosVal = 250;
                58  :   r_cosVal = 249;
                63  :   r_cosVal = 248;
                67  :   r_cosVal = 247;
                71  :   r_cosVal = 246;
                76  :   r_cosVal = 245;
                80  :   r_cosVal = 243;
                85  :   r_cosVal = 242;
                89  :   r_cosVal = 241;
                94  :   r_cosVal = 239;
                98  :   r_cosVal = 237;
                103 :   r_cosVal = 236;
                107 :   r_cosVal = 234;
                112 :   r_cosVal = 232;
                116 :   r_cosVal = 230;
                121 :   r_cosVal = 228;
                125 :   r_cosVal = 226;
                130 :   r_cosVal = 224;
                134 :   r_cosVal = 222;
                139 :   r_cosVal = 219;
                143 :   r_cosVal = 217;
                147 :   r_cosVal = 215;
                152 :   r_cosVal = 212;
                156 :   r_cosVal = 210;
                161 :   r_cosVal = 207;
                165 :   r_cosVal = 204;
                170 :   r_cosVal = 202;
                174 :   r_cosVal = 199;
                179 :   r_cosVal = 196;
                183 :   r_cosVal = 193;
                188 :   r_cosVal = 190;
                192 :   r_cosVal = 187;
                197 :   r_cosVal = 184;
                201 :   r_cosVal = 181;
                206 :   r_cosVal = 178;
                210 :   r_cosVal = 175;
                214 :   r_cosVal = 171;
                219 :   r_cosVal = 168;
                223 :   r_cosVal = 165;
                228 :   r_cosVal = 161;
                232 :   r_cosVal = 158;
                237 :   r_cosVal = 154;
                241 :   r_cosVal = 150;
                246 :   r_cosVal = 147;
                250 :   r_cosVal = 143;
                255 :   r_cosVal = 139;
                259 :   r_cosVal = 136;
                264 :   r_cosVal = 132;
                268 :   r_cosVal = 128;
                273 :   r_cosVal = 124;
                277 :   r_cosVal = 120;
                281 :   r_cosVal = 116;
                286 :   r_cosVal = 112;
                290 :   r_cosVal = 108;
                295 :   r_cosVal = 104;
                299 :   r_cosVal = 100;
                304 :   r_cosVal = 96;
                308 :   r_cosVal = 92;
                313 :   r_cosVal = 88;
                317 :   r_cosVal = 83;
                322 :   r_cosVal = 79;
                326 :   r_cosVal = 75;
                331 :   r_cosVal = 71;
                335 :   r_cosVal = 66;
                340 :   r_cosVal = 62;
                344 :   r_cosVal = 58;
                349 :   r_cosVal = 53;
                353 :   r_cosVal = 49;
                357 :   r_cosVal = 44;
                362 :   r_cosVal = 40;
                366 :   r_cosVal = 36;
                371 :   r_cosVal = 31;
                375 :   r_cosVal = 27;
                380 :   r_cosVal = 22;
                384 :   r_cosVal = 18;
                389 :   r_cosVal = 13;
                393 :   r_cosVal = 9;
                398 :   r_cosVal = 4;
                402 :   r_cosVal = 0;
                407 :   r_cosVal = -4;
                411 :   r_cosVal = -9;
                416 :   r_cosVal = -13;
                420 :   r_cosVal = -18;
                424 :   r_cosVal = -22;
                429 :   r_cosVal = -27;
                433 :   r_cosVal = -31;
                438 :   r_cosVal = -36;
                442 :   r_cosVal = -40;
                447 :   r_cosVal = -44;
                451 :   r_cosVal = -49;
                456 :   r_cosVal = -53;
                460 :   r_cosVal = -58;
                465 :   r_cosVal = -62;
                469 :   r_cosVal = -66;
                474 :   r_cosVal = -71;
                478 :   r_cosVal = -75;
                483 :   r_cosVal = -79;
                487 :   r_cosVal = -83;
                491 :   r_cosVal = -88;
                496 :   r_cosVal = -92;
                500 :   r_cosVal = -96;
                505 :   r_cosVal = -100;
                509 :   r_cosVal = -104;
                514 :   r_cosVal = -108;
                518 :   r_cosVal = -112;
                523 :   r_cosVal = -116;
                527 :   r_cosVal = -120;
                532 :   r_cosVal = -124;
                536 :   r_cosVal = -128;
                541 :   r_cosVal = -132;
                545 :   r_cosVal = -136;
                550 :   r_cosVal = -139;
                554 :   r_cosVal = -143;
                559 :   r_cosVal = -147;
                563 :   r_cosVal = -150;
                567 :   r_cosVal = -154;
                572 :   r_cosVal = -158;
                576 :   r_cosVal = -161;
                581 :   r_cosVal = -165;
                585 :   r_cosVal = -168;
                590 :   r_cosVal = -171;
                594 :   r_cosVal = -175;
                599 :   r_cosVal = -178;
                603 :   r_cosVal = -181;
                608 :   r_cosVal = -184;
                612 :   r_cosVal = -187;
                617 :   r_cosVal = -190;
                621 :   r_cosVal = -193;
                626 :   r_cosVal = -196;
                630 :   r_cosVal = -199;
                634 :   r_cosVal = -202;
                639 :   r_cosVal = -204;
                643 :   r_cosVal = -207;
                648 :   r_cosVal = -210;
                652 :   r_cosVal = -212;
                657 :   r_cosVal = -215;
                661 :   r_cosVal = -217;
                666 :   r_cosVal = -219;
                670 :   r_cosVal = -222;
                675 :   r_cosVal = -224;
                679 :   r_cosVal = -226;
                684 :   r_cosVal = -228;
                688 :   r_cosVal = -230;
                693 :   r_cosVal = -232;
                697 :   r_cosVal = -234;
                701 :   r_cosVal = -236;
                706 :   r_cosVal = -237;
                710 :   r_cosVal = -239;
                715 :   r_cosVal = -241;
                719 :   r_cosVal = -242;
                724 :   r_cosVal = -243;
                728 :   r_cosVal = -245;
                733 :   r_cosVal = -246;
                737 :   r_cosVal = -247;
                742 :   r_cosVal = -248;
                746 :   r_cosVal = -249;
                751 :   r_cosVal = -250;
                755 :   r_cosVal = -251;
                760 :   r_cosVal = -252;
                764 :   r_cosVal = -253;
                769 :   r_cosVal = -254;
                773 :   r_cosVal = -254;
                777 :   r_cosVal = -255;
                782 :   r_cosVal = -255;
                786 :   r_cosVal = -255;
                791 :   r_cosVal = -256;
                795 :   r_cosVal = -256;
                800 :   r_cosVal = -256;
                804 :   r_cosVal = -256;
            endcase
        end
    end

    assign o_cosVal_q8_8 = r_cosVal;
    
endmodule
//////////////////////////////////////////////////////////////////////////////////
module arccos_LUT (
    input       wire                                    i_reset,
    input       wire        signed      [15 : 0]        i_cosVal_q8_8,
    output      wire        signed      [15 : 0]        o_radVal_q8_8
);
                reg         signed      [15 : 0]        r_radVal;

    always @(*) begin
        if (i_reset) begin
            r_radVal = 0;
        end
        else begin
            case (i_cosVal_q8_8)
                256  : r_radVal = 0;
                256  : r_radVal = 4;
                256  : r_radVal = 9;
                256  : r_radVal = 13;
                255  : r_radVal = 18;
                255  : r_radVal = 22;
                255  : r_radVal = 27;
                254  : r_radVal = 31;
                254  : r_radVal = 36;
                253  : r_radVal = 40;
                252  : r_radVal = 45;
                251  : r_radVal = 49;
                250  : r_radVal = 54;
                249  : r_radVal = 58;
                248  : r_radVal = 63;
                247  : r_radVal = 67;
                246  : r_radVal = 71;
                245  : r_radVal = 76;
                244  : r_radVal = 78;
                243  : r_radVal = 80;
                242  : r_radVal = 85;
                241  : r_radVal = 89;
                240  : r_radVal = 92;
                239  : r_radVal = 94;
                238  : r_radVal = 96;
                237  : r_radVal = 98;
                236  : r_radVal = 103;
                235  : r_radVal = 105;
                234  : r_radVal = 107;
                233  : r_radVal = 109;
                232  : r_radVal = 112;
                231  : r_radVal = 114;
                230  : r_radVal = 116;
                229  : r_radVal = 118;
                228  : r_radVal = 121;
                227  : r_radVal = 123;
                226  : r_radVal = 125;
                225  : r_radVal = 128;
                224  : r_radVal = 130;
                223  : r_radVal = 132;
                222  : r_radVal = 134;
                221  : r_radVal = 136;
                220  : r_radVal = 137;
                219  : r_radVal = 139;
                218  : r_radVal = 140;
                217  : r_radVal = 143;
                216  : r_radVal = 145;
                215  : r_radVal = 147;
                214  : r_radVal = 149;  
                213  : r_radVal = 150;  
                212  : r_radVal = 152;
                211  : r_radVal = 154;
                210  : r_radVal = 156;
                209  : r_radVal = 158;  
                208  : r_radVal = 160;  
                207  : r_radVal = 161;
                206  : r_radVal = 163;
                205  : r_radVal = 164;  
                204  : r_radVal = 165;
                203  : r_radVal = 167;  
                202  : r_radVal = 170;
                201  : r_radVal = 172;  
                200  : r_radVal = 173;  
                199  : r_radVal = 174;
                198  : r_radVal = 176;  
                197  : r_radVal = 177;  
                196  : r_radVal = 179;
                195  : r_radVal = 181;  
                194  : r_radVal = 182;  
                193  : r_radVal = 183;
                192  : r_radVal = 185;  
                191  : r_radVal = 187;  
                190  : r_radVal = 188;
                189  : r_radVal = 190;  
                188  : r_radVal = 191;  
                187  : r_radVal = 192;
                186  : r_radVal = 194;  
                185  : r_radVal = 195;  
                184  : r_radVal = 197;
                183  : r_radVal = 199;  
                182  : r_radVal = 200;  
                181  : r_radVal = 201;
                180  : r_radVal = 203;  
                179  : r_radVal = 204;  
                178  : r_radVal = 206;
                177  : r_radVal = 208;  
                176  : r_radVal = 209;  
                175  : r_radVal = 210;
                174  : r_radVal = 212;  
                173  : r_radVal = 213;  
                172  : r_radVal = 215;  
                171  : r_radVal = 214;
                170  : r_radVal = 217;  
                169  : r_radVal = 218;  
                168  : r_radVal = 219;
                167  : r_radVal = 220;  
                166  : r_radVal = 221;  
                165  : r_radVal = 223;
                164  : r_radVal = 224;  
                163  : r_radVal = 225;
                162  : r_radVal = 227;  
                161  : r_radVal = 228;
                160  : r_radVal = 230;
                159  : r_radVal = 231;
                158  : r_radVal = 232;
                157  : r_radVal = 233;  
                156  : r_radVal = 234;  
                155  : r_radVal = 236;  
                154  : r_radVal = 237;
                153  : r_radVal = 239;  
                152  : r_radVal = 240;  
                150  : r_radVal = 241;
                149  : r_radVal = 243;  
                148  : r_radVal = 244;  
                147  : r_radVal = 246;
                146  : r_radVal = 247;  
                145  : r_radVal = 248;  
                144  : r_radVal = 249;  
                143  : r_radVal = 250;
                142  : r_radVal = 252;  
                141  : r_radVal = 253;  
                140  : r_radVal = 254;  
                139  : r_radVal = 255;
                138  : r_radVal = 257;  
                137  : r_radVal = 258;  
                136  : r_radVal = 259;
                135  : r_radVal = 261;  
                134  : r_radVal = 262;  
                133  : r_radVal = 263;  
                132  : r_radVal = 264;
                131  : r_radVal = 266;  
                130  : r_radVal = 267;  
                129  : r_radVal = 268;  
                128  : r_radVal = 268;
                127  : r_radVal = 269;  
                126  : r_radVal = 270;  
                125  : r_radVal = 270;
                124  : r_radVal = 273;
                123  : r_radVal = 274;  
                122  : r_radVal = 275;  
                121  : r_radVal = 276;  
                120  : r_radVal = 277;
                119  : r_radVal = 279;
                118  : r_radVal = 280;  
                117  : r_radVal = 281;  
                116  : r_radVal = 281;
                115  : r_radVal = 282;
                114  : r_radVal = 283;  
                113  : r_radVal = 284;
                112  : r_radVal = 286;
                111  : r_radVal = 287;  
                110  : r_radVal = 288;  
                109  : r_radVal = 289;  
                108  : r_radVal = 290;
                107  : r_radVal = 292;  
                106  : r_radVal = 293;  
                105  : r_radVal = 294;  
                104  : r_radVal = 295;
                103  : r_radVal = 297;  
                102  : r_radVal = 298;  
                101  : r_radVal = 299;  
                100  : r_radVal = 299;
                99   : r_radVal = 301;  
                98   : r_radVal = 302;  
                97   : r_radVal = 303;  
                96   : r_radVal = 304;
                95   : r_radVal = 306;  
                94   : r_radVal = 307;  
                93   : r_radVal = 308;
                92   : r_radVal = 308;
                91   : r_radVal = 310;  
                90   : r_radVal = 311;  
                89   : r_radVal = 312;  
                88   : r_radVal = 313;
                87   : r_radVal = 315;  
                86   : r_radVal = 316;  
                85   : r_radVal = 317;  
                84   : r_radVal = 318;  
                83   : r_radVal = 317;
                82   : r_radVal = 319;  
                81   : r_radVal = 320;  
                80   : r_radVal = 321;  
                79   : r_radVal = 322;
                78   : r_radVal = 323;  
                77   : r_radVal = 324;  
                76   : r_radVal = 324;
                75   : r_radVal = 326;
                74   : r_radVal = 327;  
                73   : r_radVal = 328;  
                72   : r_radVal = 329;
                71   : r_radVal = 331;
                70   : r_radVal = 332;  
                69   : r_radVal = 333;  
                68   : r_radVal = 334;  
                67   : r_radVal = 335;
                66   : r_radVal = 335;
                65   : r_radVal = 337;  
                64   : r_radVal = 338;  
                63   : r_radVal = 339;  
                62   : r_radVal = 340;
                61   : r_radVal = 341;  
                60   : r_radVal = 342;  
                59   : r_radVal = 343;  
                58   : r_radVal = 344;
                57   : r_radVal = 345;  
                56   : r_radVal = 346;  
                55   : r_radVal = 347;  
                54   : r_radVal = 348;  
                53   : r_radVal = 349;
                52   : r_radVal = 350;  
                51   : r_radVal = 351;  
                50   : r_radVal = 352;  
                49   : r_radVal = 353;
                48   : r_radVal = 354;  
                47   : r_radVal = 355;  
                46   : r_radVal = 356;  
                45   : r_radVal = 357;
                44   : r_radVal = 357;
                43   : r_radVal = 360;
                42   : r_radVal = 361;  
                41   : r_radVal = 362;  
                40   : r_radVal = 362;
                39   : r_radVal = 363;  
                38   : r_radVal = 364;  
                37   : r_radVal = 364;
                36   : r_radVal = 366;
                35   : r_radVal = 366;  
                34   : r_radVal = 367;  
                33   : r_radVal = 368;
                32   : r_radVal = 369;
                31   : r_radVal = 371;
                30   : r_radVal = 372;  
                29   : r_radVal = 373;  
                28   : r_radVal = 374;  
                27   : r_radVal = 375;
                26   : r_radVal = 376;  
                25   : r_radVal = 377;  
                24   : r_radVal = 378;  
                23   : r_radVal = 379;  
                22   : r_radVal = 380;
                21   : r_radVal = 381;  
                20   : r_radVal = 382;  
                19   : r_radVal = 383;  
                18   : r_radVal = 384;
                17   : r_radVal = 385;  
                16   : r_radVal = 386;  
                15   : r_radVal = 387;  
                14   : r_radVal = 388;  
                13   : r_radVal = 389;
                12   : r_radVal = 390;  
                11   : r_radVal = 391;  
                10   : r_radVal = 392;  
                9    : r_radVal = 393;
                8    : r_radVal = 394;  
                7    : r_radVal = 395;  
                6    : r_radVal = 395;
                5    : r_radVal = 397;  
                4    : r_radVal = 398;
                3    : r_radVal = 399;  
                2    : r_radVal = 400;  
                1    : r_radVal = 401;  
                0    : r_radVal = 402;
                -1   : r_radVal = 403;  
                -2   : r_radVal = 404;  
                -3   : r_radVal = 405;  
                -4   : r_radVal = 407;
                -5   : r_radVal = 408;  
                -6   : r_radVal = 409;
                -7   : r_radVal = 410;  
                -8   : r_radVal = 411;  
                -9   : r_radVal = 411;
                -10  : r_radVal = 412;  
                -11  : r_radVal = 413;  
                -12  : r_radVal = 414;  
                -13  : r_radVal = 416;
                -14  : r_radVal = 417;  
                -15  : r_radVal = 418;  
                -16  : r_radVal = 419;  
                -17  : r_radVal = 420;  
                -18  : r_radVal = 420;
                -19  : r_radVal = 422;  
                -20  : r_radVal = 423;  
                -21  : r_radVal = 424;
                -22  : r_radVal = 424;
                -23  : r_radVal = 426;  
                -24  : r_radVal = 427;  
                -25  : r_radVal = 428;  
                -26  : r_radVal = 429;  
                -27  : r_radVal = 429;
                -28  : r_radVal = 430;  
                -29  : r_radVal = 431;
                -30  : r_radVal = 432;  
                -31  : r_radVal = 433;
                -32  : r_radVal = 434;  
                -33  : r_radVal = 435;  
                -34  : r_radVal = 436;  
                -35  : r_radVal = 436;
                -36  : r_radVal = 438;
                -37  : r_radVal = 439;  
                -38  : r_radVal = 440;  
                -39  : r_radVal = 440;
                -40  : r_radVal = 442;
                -41  : r_radVal = 443;  
                -42  : r_radVal = 444;  
                -43  : r_radVal = 445;  
                -44  : r_radVal = 447;
                -45  : r_radVal = 448;  
                -46  : r_radVal = 449;  
                -47  : r_radVal = 450;  
                -48  : r_radVal = 451;  
                -49  : r_radVal = 451;
                -50  : r_radVal = 453;  
                -51  : r_radVal = 454;  
                -52  : r_radVal = 455;  
                -53  : r_radVal = 456;
                -54  : r_radVal = 457;  
                -55  : r_radVal = 458;  
                -56  : r_radVal = 459;  
                -57  : r_radVal = 460;  
                -58  : r_radVal = 460;
                -59  : r_radVal = 462;  
                -60  : r_radVal = 463;  
                -61  : r_radVal = 463;
                -62  : r_radVal = 465;
                -63  : r_radVal = 466;  
                -64  : r_radVal = 467;  
                -65  : r_radVal = 468;  
                -66  : r_radVal = 469;
                -67  : r_radVal = 470;
                -68  : r_radVal = 471;  
                -69  : r_radVal = 472;  
                -70  : r_radVal = 473;  
                -71  : r_radVal = 474;
                -72  : r_radVal = 476;
                -73  : r_radVal = 477;  
                -74  : r_radVal = 478;  
                -75  : r_radVal = 478;
                -76  : r_radVal = 480;  
                -77  : r_radVal = 481;  
                -78  : r_radVal = 482;  
                -79  : r_radVal = 483;
                -80  : r_radVal = 484;  
                -81  : r_radVal = 485;  
                -82  : r_radVal = 486;  
                -83  : r_radVal = 487;
                -84  : r_radVal = 488;  
                -85  : r_radVal = 489;  
                -86  : r_radVal = 490;  
                -87  : r_radVal = 491;  
                -88  : r_radVal = 491;
                -89  : r_radVal = 493;  
                -90  : r_radVal = 494;
                -91  : r_radVal = 495;  
                -92  : r_radVal = 496;
                -93  : r_radVal = 497;  
                -94  : r_radVal = 498;  
                -95  : r_radVal = 499;  
                -96  : r_radVal = 500;
                -97  : r_radVal = 501;  
                -98  : r_radVal = 502;  
                -99  : r_radVal = 503;  
                -100 : r_radVal = 505;
                -101 : r_radVal = 506;  
                -102 : r_radVal = 507;
                -103 : r_radVal = 508;  
                -104 : r_radVal = 509;
                -105 : r_radVal = 510;  
                -106 : r_radVal = 511;  
                -107 : r_radVal = 512;  
                -108 : r_radVal = 514;
                -109 : r_radVal = 515;  
                -110 : r_radVal = 516;  
                -111 : r_radVal = 517;  
                -112 : r_radVal = 518;
                -113 : r_radVal = 519;  
                -114 : r_radVal = 520;  
                -115 : r_radVal = 521;  
                -116 : r_radVal = 523;
                -117 : r_radVal = 525;
                -118 : r_radVal = 526;  
                -119 : r_radVal = 527;  
                -120 : r_radVal = 527;
                -121 : r_radVal = 528;  
                -122 : r_radVal = 529;  
                -123 : r_radVal = 531;
                -124 : r_radVal = 532;
                -125 : r_radVal = 533;  
                -126 : r_radVal = 534;  
                -127 : r_radVal = 534;
                -128 : r_radVal = 536;
                -129 : r_radVal = 537;  
                -130 : r_radVal = 538;  
                -131 : r_radVal = 539;  
                -132 : r_radVal = 541;
                -133 : r_radVal = 542;  
                -134 : r_radVal = 543;  
                -135 : r_radVal = 544;  
                -136 : r_radVal = 545;
                -137 : r_radVal = 546;  
                -138 : r_radVal = 547;  
                -139 : r_radVal = 550;
                -140 : r_radVal = 551;
                -141 : r_radVal = 552;
                -142 : r_radVal = 553;  
                -143 : r_radVal = 554;
                -144 : r_radVal = 555;  
                -145 : r_radVal = 556;  
                -146 : r_radVal = 557;  
                -147 : r_radVal = 559;
                -148 : r_radVal = 561;
                -149 : r_radVal = 562;  
                -150 : r_radVal = 563;
                -151 : r_radVal = 564;  
                -152 : r_radVal = 564;
                -153 : r_radVal = 565;
                -154 : r_radVal = 567;
                -155 : r_radVal = 568;  
                -156 : r_radVal = 569;  
                -157 : r_radVal = 570;  
                -158 : r_radVal = 572;
                -159 : r_radVal = 573;  
                -160 : r_radVal = 574;  
                -161 : r_radVal = 576;
                -162 : r_radVal = 577;  
                -163 : r_radVal = 579;
                -164 : r_radVal = 580;  
                -165 : r_radVal = 581;
                -166 : r_radVal = 582;  
                -167 : r_radVal = 583;  
                -168 : r_radVal = 585;
                -169 : r_radVal = 587;
                -170 : r_radVal = 588;  
                -171 : r_radVal = 590;
                -172 : r_radVal = 591;  
                -173 : r_radVal = 592;
                -174 : r_radVal = 593;  
                -175 : r_radVal = 594;
                -176 : r_radVal = 595;  
                -177 : r_radVal = 596;  
                -178 : r_radVal = 599;
                -179 : r_radVal = 600;  
                -180 : r_radVal = 601;  
                -181 : r_radVal = 603;
                -182 : r_radVal = 605;
                -183 : r_radVal = 606;  
                -184 : r_radVal = 608;
                -185 : r_radVal = 609;  
                -186 : r_radVal = 610;  
                -187 : r_radVal = 612;
                -188 : r_radVal = 613;  
                -189 : r_radVal = 615;
                -190 : r_radVal = 617;
                -191 : r_radVal = 618;  
                -192 : r_radVal = 619;
                -193 : r_radVal = 621;
                -194 : r_radVal = 624;
                -195 : r_radVal = 625;  
                -196 : r_radVal = 626;
                -197 : r_radVal = 628;  
                -198 : r_radVal = 629;  
                -199 : r_radVal = 630;
                -200 : r_radVal = 631;  
                -201 : r_radVal = 632;  
                -202 : r_radVal = 634;
                -203 : r_radVal = 635;  
                -204 : r_radVal = 639;
                -205 : r_radVal = 641;
                -206 : r_radVal = 642;  
                -207 : r_radVal = 643;
                -208 : r_radVal = 644;  
                -209 : r_radVal = 646;
                -210 : r_radVal = 648;
                -211 : r_radVal = 650;
                -212 : r_radVal = 652;
                -213 : r_radVal = 654;
                -214 : r_radVal = 656;
                -215 : r_radVal = 658;
                -216 : r_radVal = 660;
                -217 : r_radVal = 662;
                -218 : r_radVal = 664;
                -219 : r_radVal = 666;
                -220 : r_radVal = 668;  
                -221 : r_radVal = 669;  
                -222 : r_radVal = 670;
                -223 : r_radVal = 673;
                -224 : r_radVal = 675;
                -225 : r_radVal = 677;  
                -226 : r_radVal = 679;
                -227 : r_radVal = 681;  
                -228 : r_radVal = 684;
                -229 : r_radVal = 686;  
                -230 : r_radVal = 688;
                -231 : r_radVal = 690;
                -232 : r_radVal = 693;
                -233 : r_radVal = 695;  
                -234 : r_radVal = 697;
                -235 : r_radVal = 699;
                -236 : r_radVal = 701;
                -237 : r_radVal = 706;
                -238 : r_radVal = 708;  
                -239 : r_radVal = 710;
                -240 : r_radVal = 712;
                -241 : r_radVal = 715;
                -242 : r_radVal = 719;
                -243 : r_radVal = 724;
                -244 : r_radVal = 726;
                -245 : r_radVal = 728;
                -246 : r_radVal = 733;
                -247 : r_radVal = 737;
                -248 : r_radVal = 742;
                -249 : r_radVal = 746;
                -250 : r_radVal = 751;
                -251 : r_radVal = 755;
                -252 : r_radVal = 760;
                -253 : r_radVal = 764;
                -254 : r_radVal = 769;
                -255 : r_radVal = 777;
                -256 : r_radVal = 791;
                default : r_radVal = r_radVal;
            endcase
        end
    end

    assign o_radVal_q8_8 = r_radVal;
endmodule
//////////////////////////////////////////////////////////////////////////////////
module arctan_LUT (
    input       wire                                    i_reset,
    input       wire        signed      [15 : 0]        i_tanVal_q8_8,
    output      wire        signed      [15 : 0]        o_radVal_q8_8
);
                reg         signed      [15 : 0]        r_radVal;

    always @(*) begin
        if (i_reset) begin
            r_radVal = 0;
        end
        else begin
            case (i_tanVal_q8_8)
                0       :   r_radVal = 0;
                256     :   r_radVal = 201;
                128     :   r_radVal = 119;
                85      :   r_radVal = 82;
                64      :   r_radVal = 63;
                51      :   r_radVal = 51;
                43      :   r_radVal = 42;
                37      :   r_radVal = 36;
                32      :   r_radVal = 32;
                28      :   r_radVal = 28;
                26      :   r_radVal = 26;
                23      :   r_radVal = 23;
                21      :   r_radVal = 21;
                20      :   r_radVal = 20;
                18      :   r_radVal = 18;
                17      :   r_radVal = 17;
                16      :   r_radVal = 16;
                15      :   r_radVal = 15;
                14      :   r_radVal = 14;
                13      :   r_radVal = 13;
                13      :   r_radVal = 13;
                512     :   r_radVal = 283;
                256     :   r_radVal = 201;
                171     :   r_radVal = 151;
                128     :   r_radVal = 119;
                102     :   r_radVal = 97;
                85      :   r_radVal = 82;
                73      :   r_radVal = 71;
                64      :   r_radVal = 63;
                57      :   r_radVal = 56;
                51      :   r_radVal = 51;
                47      :   r_radVal = 46;
                43      :   r_radVal = 42;
                39      :   r_radVal = 39;
                37      :   r_radVal = 36;
                34      :   r_radVal = 34;
                32      :   r_radVal = 32;
                30      :   r_radVal = 30;
                28      :   r_radVal = 28;
                27      :   r_radVal = 27;
                26      :   r_radVal = 26;
                768     :   r_radVal = 320;
                384     :   r_radVal = 252;
                256     :   r_radVal = 201;
                192     :   r_radVal = 165;
                154     :   r_radVal = 138;
                128     :   r_radVal = 119;
                110     :   r_radVal = 104;
                96      :   r_radVal = 92;
                85      :   r_radVal = 82;
                77      :   r_radVal = 75;
                70      :   r_radVal = 68;
                64      :   r_radVal = 63;
                59      :   r_radVal = 58;
                55      :   r_radVal = 54;
                51      :   r_radVal = 51;
                48      :   r_radVal = 47;
                45      :   r_radVal = 45;
                43      :   r_radVal = 42;
                40      :   r_radVal = 40;
                38      :   r_radVal = 38;
                1024    :   r_radVal = 339;
                512     :   r_radVal = 283;
                341     :   r_radVal = 237;
                256     :   r_radVal = 201;
                205     :   r_radVal = 173;
                171     :   r_radVal = 151;
                146     :   r_radVal = 133;
                128     :   r_radVal = 119;
                114     :   r_radVal = 107;
                102     :   r_radVal = 97;
                93      :   r_radVal = 89;
                85      :   r_radVal = 82;
                79      :   r_radVal = 76;
                73      :   r_radVal = 71;
                68      :   r_radVal = 67;
                64      :   r_radVal = 63;
                60      :   r_radVal = 59;
                57      :   r_radVal = 56;
                54      :   r_radVal = 53;
                51      :   r_radVal = 51;
                1280    :   r_radVal = 352;
                640     :   r_radVal = 305;
                427     :   r_radVal = 264;
                320     :   r_radVal = 229;
                256     :   r_radVal = 201;
                213     :   r_radVal = 178;
                183     :   r_radVal = 159;
                160     :   r_radVal = 143;
                142     :   r_radVal = 130;
                128     :   r_radVal = 119;
                116     :   r_radVal = 109;
                107     :   r_radVal = 101;
                98      :   r_radVal = 94;
                91      :   r_radVal = 88;
                85      :   r_radVal = 82;
                80      :   r_radVal = 78;
                75      :   r_radVal = 73;
                71      :   r_radVal = 69;
                67      :   r_radVal = 66;
                64      :   r_radVal = 63;
                1536    :   r_radVal = 360;
                768     :   r_radVal = 320;
                512     :   r_radVal = 283;
                384     :   r_radVal = 252;
                307     :   r_radVal = 224;
                256     :   r_radVal = 201;
                219     :   r_radVal = 181;
                192     :   r_radVal = 165;
                171     :   r_radVal = 151;
                154     :   r_radVal = 138;
                140     :   r_radVal = 128;
                128     :   r_radVal = 119;
                118     :   r_radVal = 111;
                110     :   r_radVal = 104;
                102     :   r_radVal = 97;
                96      :   r_radVal = 92;
                90      :   r_radVal = 87;
                85      :   r_radVal = 82;
                81      :   r_radVal = 78;
                77      :   r_radVal = 75;
                1792    :   r_radVal = 366;
                896     :   r_radVal = 331;
                597     :   r_radVal = 298;
                448     :   r_radVal = 269;
                358     :   r_radVal = 243;
                299     :   r_radVal = 221;
                256     :   r_radVal = 201;
                224     :   r_radVal = 184;
                199     :   r_radVal = 169;
                179     :   r_radVal = 156;
                163     :   r_radVal = 145;
                149     :   r_radVal = 135;
                138     :   r_radVal = 126;
                128     :   r_radVal = 119;
                119     :   r_radVal = 112;
                112     :   r_radVal = 106;
                105     :   r_radVal = 100;
                100     :   r_radVal = 95;
                94      :   r_radVal = 90;
                90      :   r_radVal = 86;
                2048    :   r_radVal = 370;
                1024    :   r_radVal = 339;
                683     :   r_radVal = 310;
                512     :   r_radVal = 283;
                410     :   r_radVal = 259;
                341     :   r_radVal = 237;
                293     :   r_radVal = 218;
                256     :   r_radVal = 201;
                228     :   r_radVal = 186;
                205     :   r_radVal = 173;
                186     :   r_radVal = 161;
                171     :   r_radVal = 151;
                158     :   r_radVal = 141;
                146     :   r_radVal = 133;
                137     :   r_radVal = 125;
                128     :   r_radVal = 119;
                120     :   r_radVal = 113;
                114     :   r_radVal = 107;
                108     :   r_radVal = 102;
                102     :   r_radVal = 97;
                2304    :   r_radVal = 374;
                1152    :   r_radVal = 346;
                768     :   r_radVal = 320;
                576     :   r_radVal = 295;
                461     :   r_radVal = 272;
                384     :   r_radVal = 252;
                329     :   r_radVal = 233;
                288     :   r_radVal = 216;
                256     :   r_radVal = 201;
                230     :   r_radVal = 188;
                209     :   r_radVal = 176;
                192     :   r_radVal = 165;
                177     :   r_radVal = 155;
                165     :   r_radVal = 146;
                154     :   r_radVal = 138;
                144     :   r_radVal = 131;
                136     :   r_radVal = 125;
                128     :   r_radVal = 119;
                121     :   r_radVal = 113;
                115     :   r_radVal = 108;
                2560    :   r_radVal = 377;
                1280    :   r_radVal = 352;
                853     :   r_radVal = 328;
                640     :   r_radVal = 305;
                512     :   r_radVal = 283;
                427     :   r_radVal = 264;
                366     :   r_radVal = 246;
                320     :   r_radVal = 229;
                284     :   r_radVal = 215;
                256     :   r_radVal = 201;
                233     :   r_radVal = 189;
                213     :   r_radVal = 178;
                197     :   r_radVal = 168;
                183     :   r_radVal = 159;
                171     :   r_radVal = 151;
                160     :   r_radVal = 143;
                151     :   r_radVal = 136;
                142     :   r_radVal = 130;
                135     :   r_radVal = 124;
                128     :   r_radVal = 119;
                2816    :   r_radVal = 379;
                1408    :   r_radVal = 356;
                939     :   r_radVal = 334;
                704     :   r_radVal = 313;
                563     :   r_radVal = 293;
                469     :   r_radVal = 274;
                402     :   r_radVal = 257;
                352     :   r_radVal = 241;
                313     :   r_radVal = 227;
                282     :   r_radVal = 213;
                256     :   r_radVal = 201;
                235     :   r_radVal = 190;
                217     :   r_radVal = 180;
                201     :   r_radVal = 170;
                188     :   r_radVal = 162;
                176     :   r_radVal = 154;
                166     :   r_radVal = 147;
                156     :   r_radVal = 140;
                148     :   r_radVal = 134;
                141     :   r_radVal = 129;
                3072    :   r_radVal = 381;
                1536    :   r_radVal = 360;
                1024    :   r_radVal = 339;
                768     :   r_radVal = 320;
                614     :   r_radVal = 301;
                512     :   r_radVal = 283;
                439     :   r_radVal = 267;
                384     :   r_radVal = 252;
                341     :   r_radVal = 237;
                307     :   r_radVal = 224;
                279     :   r_radVal = 212;
                256     :   r_radVal = 201;
                236     :   r_radVal = 191;
                219     :   r_radVal = 181;
                205     :   r_radVal = 173;
                192     :   r_radVal = 165;
                181     :   r_radVal = 157;
                171     :   r_radVal = 151;
                162     :   r_radVal = 144;
                154     :   r_radVal = 138;
                3328    :   r_radVal = 382;
                1664    :   r_radVal = 363;
                1109    :   r_radVal = 344;
                832     :   r_radVal = 326;
                666     :   r_radVal = 308;
                555     :   r_radVal = 291;
                475     :   r_radVal = 276;
                416     :   r_radVal = 261;
                370     :   r_radVal = 247;
                333     :   r_radVal = 234;
                303     :   r_radVal = 222;
                277     :   r_radVal = 211;
                256     :   r_radVal = 201;
                238     :   r_radVal = 192;
                222     :   r_radVal = 183;
                208     :   r_radVal = 175;
                196     :   r_radVal = 167;
                185     :   r_radVal = 160;
                175     :   r_radVal = 154;
                166     :   r_radVal = 148;
                3584    :   r_radVal = 384;
                1792    :   r_radVal = 366;
                1195    :   r_radVal = 348;
                896     :   r_radVal = 331;
                717     :   r_radVal = 314;
                597     :   r_radVal = 298;
                512     :   r_radVal = 283;
                448     :   r_radVal = 269;
                398     :   r_radVal = 256;
                358     :   r_radVal = 243;
                326     :   r_radVal = 232;
                299     :   r_radVal = 221;
                276     :   r_radVal = 211;
                256     :   r_radVal = 201;
                239     :   r_radVal = 192;
                224     :   r_radVal = 184;
                211     :   r_radVal = 176;
                199     :   r_radVal = 169;
                189     :   r_radVal = 163;
                179     :   r_radVal = 156;
                3840    :   r_radVal = 385;
                1920    :   r_radVal = 368;
                1280    :   r_radVal = 352;
                960     :   r_radVal = 335;
                768     :   r_radVal = 320;
                640     :   r_radVal = 305;
                549     :   r_radVal = 290;
                480     :   r_radVal = 277;
                427     :   r_radVal = 264;
                384     :   r_radVal = 252;
                349     :   r_radVal = 240;
                320     :   r_radVal = 229;
                295     :   r_radVal = 219;
                274     :   r_radVal = 210;
                256     :   r_radVal = 201;
                240     :   r_radVal = 193;
                226     :   r_radVal = 185;
                213     :   r_radVal = 178;
                202     :   r_radVal = 171;
                192     :   r_radVal = 165;
                4096    :   r_radVal = 386;
                2048    :   r_radVal = 370;
                1365    :   r_radVal = 355;
                1024    :   r_radVal = 339;
                819     :   r_radVal = 325;
                683     :   r_radVal = 310;
                585     :   r_radVal = 297;
                512     :   r_radVal = 283;
                455     :   r_radVal = 271;
                410     :   r_radVal = 259;
                372     :   r_radVal = 248;
                341     :   r_radVal = 237;
                315     :   r_radVal = 227;
                293     :   r_radVal = 218;
                273     :   r_radVal = 209;
                256     :   r_radVal = 201;
                241     :   r_radVal = 193;
                228     :   r_radVal = 186;
                216     :   r_radVal = 179;
                205     :   r_radVal = 173;
                4352    :   r_radVal = 387;
                2176    :   r_radVal = 372;
                1451    :   r_radVal = 357;
                1088    :   r_radVal = 343;
                870     :   r_radVal = 329;
                725     :   r_radVal = 315;
                622     :   r_radVal = 302;
                544     :   r_radVal = 290;
                484     :   r_radVal = 277;
                435     :   r_radVal = 266;
                396     :   r_radVal = 255;
                363     :   r_radVal = 245;
                335     :   r_radVal = 235;
                311     :   r_radVal = 226;
                290     :   r_radVal = 217;
                272     :   r_radVal = 209;
                256     :   r_radVal = 201;
                242     :   r_radVal = 194;
                229     :   r_radVal = 187;
                218     :   r_radVal = 180;
                4608    :   r_radVal = 388;
                2304    :   r_radVal = 374;
                1536    :   r_radVal = 360;
                1152    :   r_radVal = 346;
                922     :   r_radVal = 333;
                768     :   r_radVal = 320;
                658     :   r_radVal = 307;
                576     :   r_radVal = 295;
                512     :   r_radVal = 283;
                461     :   r_radVal = 272;
                419     :   r_radVal = 262;
                384     :   r_radVal = 252;
                354     :   r_radVal = 242;
                329     :   r_radVal = 233;
                307     :   r_radVal = 224;
                288     :   r_radVal = 216;
                271     :   r_radVal = 208;
                256     :   r_radVal = 201;
                243     :   r_radVal = 194;
                230     :   r_radVal = 188;
                4864    :   r_radVal = 389;
                2432    :   r_radVal = 375;
                1621    :   r_radVal = 362;
                1216    :   r_radVal = 349;
                973     :   r_radVal = 336;
                811     :   r_radVal = 324;
                695     :   r_radVal = 312;
                608     :   r_radVal = 300;
                540     :   r_radVal = 289;
                486     :   r_radVal = 278;
                442     :   r_radVal = 268;
                405     :   r_radVal = 258;
                374     :   r_radVal = 249;
                347     :   r_radVal = 240;
                324     :   r_radVal = 231;
                304     :   r_radVal = 223;
                286     :   r_radVal = 215;
                270     :   r_radVal = 208;
                256     :   r_radVal = 201;
                243     :   r_radVal = 194;
                6912    :   r_radVal = 393;
                2508    :   r_radVal = 376;
                1745    :   r_radVal = 365;
                1280    :   r_radVal = 352;
                992     :   r_radVal = 337;
                818     :   r_radVal = 324;
                685     :   r_radVal = 311;
                591     :   r_radVal = 297;
                509     :   r_radVal = 283;
                444     :   r_radVal = 268;
                390     :   r_radVal = 253;
                340     :   r_radVal = 237;
                299     :   r_radVal = 221;
                262     :   r_radVal = 204;
                225     :   r_radVal = 185;
                192     :   r_radVal = 165;
                158     :   r_radVal = 142;
                124     :   r_radVal = 115;
                84      :   r_radVal = 81;
                6912    :   r_radVal = 393;
                4480    :   r_radVal = 388;
                2261    :   r_radVal = 373;
                1642    :   r_radVal = 363;
                1243    :   r_radVal = 350;
                969     :   r_radVal = 336;
                811     :   r_radVal = 324;
                676     :   r_radVal = 309;
                582     :   r_radVal = 296;
                507     :   r_radVal = 282;
                442     :   r_radVal = 268;
                387     :   r_radVal = 253;
                340     :   r_radVal = 237;
                298     :   r_radVal = 220;
                260     :   r_radVal = 203;
                224     :   r_radVal = 184;
                192     :   r_radVal = 165;
                157     :   r_radVal = 141;
                123     :   r_radVal = 115;
                82      :   r_radVal = 79;
                2508    :   r_radVal = 376;
                2261    :   r_radVal = 373;
                1792    :   r_radVal = 366;
                1456    :   r_radVal = 358;
                1136    :   r_radVal = 345;
                913     :   r_radVal = 332;
                762     :   r_radVal = 319;
                661     :   r_radVal = 308;
                564     :   r_radVal = 293;
                493     :   r_radVal = 280;
                433     :   r_radVal = 265;
                380     :   r_radVal = 250;
                334     :   r_radVal = 235;
                294     :   r_radVal = 219;
                256     :   r_radVal = 201;
                221     :   r_radVal = 182;
                188     :   r_radVal = 162;
                154     :   r_radVal = 139;
                120     :   r_radVal = 112;
                79      :   r_radVal = 77;
                1745    :   r_radVal = 365;
                1642    :   r_radVal = 363;
                1456    :   r_radVal = 358;
                1179    :   r_radVal = 347;
                992     :   r_radVal = 337;
                839     :   r_radVal = 326;
                723     :   r_radVal = 315;
                622     :   r_radVal = 302;
                545     :   r_radVal = 290;
                476     :   r_radVal = 276;
                418     :   r_radVal = 261;
                370     :   r_radVal = 247;
                325     :   r_radVal = 231;
                286     :   r_radVal = 215;
                250     :   r_radVal = 198;
                216     :   r_radVal = 179;
                182     :   r_radVal = 158;
                149     :   r_radVal = 135;
                115     :   r_radVal = 108;
                73      :   r_radVal = 71;
                1280    :   r_radVal = 352;
                1243    :   r_radVal = 350;
                1136    :   r_radVal = 345;
                992     :   r_radVal = 337;
                876     :   r_radVal = 329;
                758     :   r_radVal = 319;
                663     :   r_radVal = 308;
                582     :   r_radVal = 296;
                512     :   r_radVal = 283;
                454     :   r_radVal = 271;
                401     :   r_radVal = 257;
                355     :   r_radVal = 242;
                313     :   r_radVal = 227;
                276     :   r_radVal = 211;
                241     :   r_radVal = 193;
                208     :   r_radVal = 175;
                175     :   r_radVal = 154;
                143     :   r_radVal = 130;
                107     :   r_radVal = 101;
                63      :   r_radVal = 62;
                992     :   r_radVal = 337;
                969     :   r_radVal = 336;
                913     :   r_radVal = 332;
                839     :   r_radVal = 326;
                758     :   r_radVal = 319;
                676     :   r_radVal = 309;
                603     :   r_radVal = 299;
                541     :   r_radVal = 289;
                480     :   r_radVal = 277;
                428     :   r_radVal = 264;
                380     :   r_radVal = 250;
                338     :   r_radVal = 236;
                299     :   r_radVal = 221;
                264     :   r_radVal = 205;
                231     :   r_radVal = 188;
                198     :   r_radVal = 169;
                167     :   r_radVal = 148;
                134     :   r_radVal = 123;
                98      :   r_radVal = 94;
                48      :   r_radVal = 47;
                818     :   r_radVal = 324;
                811     :   r_radVal = 324;
                762     :   r_radVal = 319;
                723     :   r_radVal = 315;
                663     :   r_radVal = 308;
                603     :   r_radVal = 299;
                548     :   r_radVal = 290;
                493     :   r_radVal = 280;
                444     :   r_radVal = 268;
                400     :   r_radVal = 256;
                356     :   r_radVal = 243;
                318     :   r_radVal = 229;
                283     :   r_radVal = 214;
                250     :   r_radVal = 198;
                218     :   r_radVal = 181;
                187     :   r_radVal = 162;
                156     :   r_radVal = 140;
                123     :   r_radVal = 115;
                85      :   r_radVal = 82;
                22      :   r_radVal = 22;
                685     :   r_radVal = 311;
                676     :   r_radVal = 309;
                661     :   r_radVal = 308;
                622     :   r_radVal = 302;
                582     :   r_radVal = 296;
                541     :   r_radVal = 289;
                493     :   r_radVal = 280;
                452     :   r_radVal = 270;
                408     :   r_radVal = 259;
                370     :   r_radVal = 247;
                332     :   r_radVal = 234;
                298     :   r_radVal = 220;
                265     :   r_radVal = 205;
                233     :   r_radVal = 189;
                203     :   r_radVal = 172;
                174     :   r_radVal = 153;
                143     :   r_radVal = 130;
                110     :   r_radVal = 104;
                69      :   r_radVal = 67;
                591     :   r_radVal = 297;
                582     :   r_radVal = 296;
                564     :   r_radVal = 293;
                545     :   r_radVal = 290;
                512     :   r_radVal = 283;
                480     :   r_radVal = 277;
                444     :   r_radVal = 268;
                408     :   r_radVal = 259;
                375     :   r_radVal = 249;
                340     :   r_radVal = 237;
                307     :   r_radVal = 224;
                276     :   r_radVal = 211;
                246     :   r_radVal = 196;
                217     :   r_radVal = 180;
                188     :   r_radVal = 162;
                158     :   r_radVal = 142;
                128     :   r_radVal = 119;
                94      :   r_radVal = 90;
                46      :   r_radVal = 46;
                509     :   r_radVal = 283;
                507     :   r_radVal = 282;
                493     :   r_radVal = 280;
                476     :   r_radVal = 276;
                454     :   r_radVal = 271;
                428     :   r_radVal = 264;
                400     :   r_radVal = 256;
                370     :   r_radVal = 247;
                340     :   r_radVal = 237;
                310     :   r_radVal = 225;
                282     :   r_radVal = 213;
                254     :   r_radVal = 200;
                225     :   r_radVal = 185;
                198     :   r_radVal = 169;
                170     :   r_radVal = 150;
                142     :   r_radVal = 130;
                111     :   r_radVal = 105;
                73      :   r_radVal = 71;
                444     :   r_radVal = 268;
                442     :   r_radVal = 268;
                433     :   r_radVal = 265;
                418     :   r_radVal = 261;
                401     :   r_radVal = 257;
                380     :   r_radVal = 250;
                356     :   r_radVal = 243;
                332     :   r_radVal = 234;
                307     :   r_radVal = 224;
                282     :   r_radVal = 213;
                256     :   r_radVal = 201;
                231     :   r_radVal = 188;
                205     :   r_radVal = 173;
                179     :   r_radVal = 156;
                152     :   r_radVal = 137;
                123     :   r_radVal = 115;
                90      :   r_radVal = 87;
                45      :   r_radVal = 45;
                390     :   r_radVal = 253;
                387     :   r_radVal = 253;
                380     :   r_radVal = 250;
                370     :   r_radVal = 247;
                355     :   r_radVal = 242;
                338     :   r_radVal = 236;
                318     :   r_radVal = 229;
                298     :   r_radVal = 220;
                276     :   r_radVal = 211;
                254     :   r_radVal = 200;
                231     :   r_radVal = 188;
                207     :   r_radVal = 174;
                182     :   r_radVal = 158;
                157     :   r_radVal = 141;
                131     :   r_radVal = 121;
                101     :   r_radVal = 96;
                63      :   r_radVal = 62;
                340     :   r_radVal = 237;
                340     :   r_radVal = 237;
                334     :   r_radVal = 235;
                325     :   r_radVal = 231;
                313     :   r_radVal = 227;
                299     :   r_radVal = 221;
                283     :   r_radVal = 214;
                265     :   r_radVal = 205;
                246     :   r_radVal = 196;
                225     :   r_radVal = 185;
                205     :   r_radVal = 173;
                182     :   r_radVal = 158;
                160     :   r_radVal = 143;
                135     :   r_radVal = 124;
                107     :   r_radVal = 101;
                74      :   r_radVal = 72;
                299     :   r_radVal = 221;
                298     :   r_radVal = 220;
                294     :   r_radVal = 219;
                286     :   r_radVal = 215;
                276     :   r_radVal = 211;
                264     :   r_radVal = 205;
                250     :   r_radVal = 198;
                233     :   r_radVal = 189;
                217     :   r_radVal = 180;
                198     :   r_radVal = 169;
                179     :   r_radVal = 156;
                157     :   r_radVal = 141;
                135     :   r_radVal = 124;
                110     :   r_radVal = 104;
                79      :   r_radVal = 77;
                31      :   r_radVal = 31;
                262     :   r_radVal = 204;
                260     :   r_radVal = 203;
                256     :   r_radVal = 201;
                250     :   r_radVal = 198;
                241     :   r_radVal = 193;
                231     :   r_radVal = 188;
                218     :   r_radVal = 181;
                203     :   r_radVal = 172;
                188     :   r_radVal = 162;
                170     :   r_radVal = 150;
                152     :   r_radVal = 137;
                131     :   r_radVal = 121;
                107     :   r_radVal = 101;
                79      :   r_radVal = 77;
                38      :   r_radVal = 38;
                225     :   r_radVal = 185;
                224     :   r_radVal = 184;
                221     :   r_radVal = 182;
                216     :   r_radVal = 179;
                208     :   r_radVal = 175;
                198     :   r_radVal = 169;
                187     :   r_radVal = 162;
                174     :   r_radVal = 153;
                158     :   r_radVal = 142;
                142     :   r_radVal = 130;
                123     :   r_radVal = 115;
                101     :   r_radVal = 96;
                74      :   r_radVal = 72;
                31      :   r_radVal = 31;
                192     :   r_radVal = 165;
                192     :   r_radVal = 165;
                188     :   r_radVal = 162;
                182     :   r_radVal = 158;
                175     :   r_radVal = 154;
                167     :   r_radVal = 148;
                156     :   r_radVal = 140;
                143     :   r_radVal = 130;
                128     :   r_radVal = 119;
                111     :   r_radVal = 105;
                90      :   r_radVal = 87;
                63      :   r_radVal = 62;
                158     :   r_radVal = 142;
                157     :   r_radVal = 141;
                154     :   r_radVal = 139;
                149     :   r_radVal = 135;
                143     :   r_radVal = 130;
                134     :   r_radVal = 123;
                123     :   r_radVal = 115;
                110     :   r_radVal = 104;
                94      :   r_radVal = 90;
                73      :   r_radVal = 71;
                45      :   r_radVal = 45;
                124     :   r_radVal = 115;
                123     :   r_radVal = 115;
                120     :   r_radVal = 112;
                115     :   r_radVal = 108;
                107     :   r_radVal = 101;
                98      :   r_radVal = 94;
                85      :   r_radVal = 82;
                69      :   r_radVal = 67;
                46      :   r_radVal = 46;
                84      :   r_radVal = 81;
                82      :   r_radVal = 79;
                79      :   r_radVal = 77;
                73      :   r_radVal = 71;
                63      :   r_radVal = 62;
                48      :   r_radVal = 47;
                22      :   r_radVal = 22;
                256     :   r_radVal = 201;
                128     :   r_radVal = 119;
                85      :   r_radVal = 82;
                64      :   r_radVal = 63;
                51      :   r_radVal = 50;
                42      :   r_radVal = 42;
                36      :   r_radVal = 36;
                32      :   r_radVal = 32;
                28      :   r_radVal = 28;
                25      :   r_radVal = 25;
                23      :   r_radVal = 23;
                21      :   r_radVal = 21;
                19      :   r_radVal = 19;
                18      :   r_radVal = 18;
                17      :   r_radVal = 17;
                16      :   r_radVal = 16;
                15      :   r_radVal = 15;
                14      :   r_radVal = 14;
                13      :   r_radVal = 13;
                0       :   r_radVal = 0;
                512     :   r_radVal = 283;
                256     :   r_radVal = 201;
                170     :   r_radVal = 150;
                128     :   r_radVal = 119;
                102     :   r_radVal = 97;
                85      :   r_radVal = 82;
                73      :   r_radVal = 71;
                64      :   r_radVal = 63;
                56      :   r_radVal = 55;
                51      :   r_radVal = 50;
                46      :   r_radVal = 46;
                42      :   r_radVal = 42;
                39      :   r_radVal = 39;
                36      :   r_radVal = 36;
                34      :   r_radVal = 34;
                32      :   r_radVal = 32;
                30      :   r_radVal = 30;
                28      :   r_radVal = 28;
                26      :   r_radVal = 26;
                0       :   r_radVal = 0;
                768     :   r_radVal = 320;
                384     :   r_radVal = 252;
                256     :   r_radVal = 201;
                192     :   r_radVal = 165;
                153     :   r_radVal = 138;
                128     :   r_radVal = 119;
                109     :   r_radVal = 103;
                96      :   r_radVal = 92;
                85      :   r_radVal = 82;
                76      :   r_radVal = 74;
                69      :   r_radVal = 67;
                64      :   r_radVal = 63;
                59      :   r_radVal = 58;
                54      :   r_radVal = 53;
                51      :   r_radVal = 50;
                48      :   r_radVal = 47;
                45      :   r_radVal = 45;
                42      :   r_radVal = 42;
                40      :   r_radVal = 40;
                0       :   r_radVal = 0;
                1024    :   r_radVal = 339;
                512     :   r_radVal = 283;
                341     :   r_radVal = 237;
                256     :   r_radVal = 201;
                204     :   r_radVal = 172;
                170     :   r_radVal = 150;
                146     :   r_radVal = 133;
                128     :   r_radVal = 119;
                113     :   r_radVal = 106;
                102     :   r_radVal = 97;
                93      :   r_radVal = 89;
                85      :   r_radVal = 82;
                78      :   r_radVal = 76;
                73      :   r_radVal = 71;
                68      :   r_radVal = 66;
                64      :   r_radVal = 63;
                60      :   r_radVal = 59;
                56      :   r_radVal = 55;
                53      :   r_radVal = 52;
                0       :   r_radVal = 0;
                1280    :   r_radVal = 352;
                640     :   r_radVal = 305;
                426     :   r_radVal = 264;
                320     :   r_radVal = 229;
                256     :   r_radVal = 201;
                213     :   r_radVal = 178;
                182     :   r_radVal = 158;
                160     :   r_radVal = 143;
                142     :   r_radVal = 130;
                128     :   r_radVal = 119;
                116     :   r_radVal = 109;
                106     :   r_radVal = 100;
                98      :   r_radVal = 94;
                91      :   r_radVal = 87;
                85      :   r_radVal = 82;
                80      :   r_radVal = 78;
                75      :   r_radVal = 73;
                71      :   r_radVal = 69;
                67      :   r_radVal = 66;
                0       :   r_radVal = 0;
                1536    :   r_radVal = 360;
                768     :   r_radVal = 320;
                512     :   r_radVal = 283;
                384     :   r_radVal = 252;
                307     :   r_radVal = 224;
                256     :   r_radVal = 201;
                219     :   r_radVal = 181;
                192     :   r_radVal = 165;
                170     :   r_radVal = 150;
                153     :   r_radVal = 138;
                139     :   r_radVal = 127;
                128     :   r_radVal = 119;
                118     :   r_radVal = 111;
                109     :   r_radVal = 103;
                102     :   r_radVal = 97;
                96      :   r_radVal = 92;
                90      :   r_radVal = 87;
                85      :   r_radVal = 82;
                80      :   r_radVal = 78;
                0       :   r_radVal = 0;
                1792    :   r_radVal = 366;
                896     :   r_radVal = 331;
                597     :   r_radVal = 298;
                448     :   r_radVal = 269;
                358     :   r_radVal = 243;
                298     :   r_radVal = 220;
                256     :   r_radVal = 201;
                224     :   r_radVal = 184;
                199     :   r_radVal = 169;
                179     :   r_radVal = 156;
                162     :   r_radVal = 144;
                149     :   r_radVal = 135;
                137     :   r_radVal = 126;
                128     :   r_radVal = 119;
                119     :   r_radVal = 111;
                112     :   r_radVal = 106;
                105     :   r_radVal = 100;
                99      :   r_radVal = 94;
                0       :   r_radVal = 0;
                2048    :   r_radVal = 370;
                1024    :   r_radVal = 339;
                682     :   r_radVal = 310;
                512     :   r_radVal = 283;
                409     :   r_radVal = 259;
                341     :   r_radVal = 237;
                292     :   r_radVal = 218;
                256     :   r_radVal = 201;
                227     :   r_radVal = 186;
                204     :   r_radVal = 172;
                186     :   r_radVal = 161;
                170     :   r_radVal = 150;
                157     :   r_radVal = 141;
                146     :   r_radVal = 133;
                136     :   r_radVal = 125;
                128     :   r_radVal = 119;
                120     :   r_radVal = 112;
                113     :   r_radVal = 106;
                0       :   r_radVal = 0;
                2304    :   r_radVal = 374;
                1152    :   r_radVal = 346;
                768     :   r_radVal = 320;
                576     :   r_radVal = 295;
                460     :   r_radVal = 272;
                384     :   r_radVal = 252;
                329     :   r_radVal = 233;
                288     :   r_radVal = 216;
                256     :   r_radVal = 201;
                230     :   r_radVal = 187;
                209     :   r_radVal = 175;
                192     :   r_radVal = 165;
                177     :   r_radVal = 155;
                164     :   r_radVal = 146;
                153     :   r_radVal = 138;
                144     :   r_radVal = 131;
                135     :   r_radVal = 124;
                0       :   r_radVal = 0;
                2560    :   r_radVal = 377;
                1280    :   r_radVal = 352;
                853     :   r_radVal = 327;
                640     :   r_radVal = 305;
                512     :   r_radVal = 283;
                426     :   r_radVal = 264;
                365     :   r_radVal = 246;
                320     :   r_radVal = 229;
                284     :   r_radVal = 214;
                256     :   r_radVal = 201;
                232     :   r_radVal = 188;
                213     :   r_radVal = 178;
                196     :   r_radVal = 167;
                182     :   r_radVal = 158;
                170     :   r_radVal = 150;
                160     :   r_radVal = 143;
                150     :   r_radVal = 136;
                0       :   r_radVal = 0;
                2816    :   r_radVal = 379;
                1408    :   r_radVal = 356;
                938     :   r_radVal = 334;
                704     :   r_radVal = 313;
                563     :   r_radVal = 293;
                469     :   r_radVal = 274;
                402     :   r_radVal = 257;
                352     :   r_radVal = 241;
                312     :   r_radVal = 226;
                281     :   r_radVal = 213;
                256     :   r_radVal = 201;
                234     :   r_radVal = 190;
                216     :   r_radVal = 179;
                201     :   r_radVal = 170;
                187     :   r_radVal = 162;
                176     :   r_radVal = 154;
                0       :   r_radVal = 0;
                3072    :   r_radVal = 381;
                1536    :   r_radVal = 360;
                1024    :   r_radVal = 339;
                768     :   r_radVal = 320;
                614     :   r_radVal = 301;
                512     :   r_radVal = 283;
                438     :   r_radVal = 267;
                384     :   r_radVal = 252;
                341     :   r_radVal = 237;
                307     :   r_radVal = 224;
                279     :   r_radVal = 212;
                256     :   r_radVal = 201;
                236     :   r_radVal = 191;
                219     :   r_radVal = 181;
                204     :   r_radVal = 172;
                0       :   r_radVal = 0;
                3328    :   r_radVal = 382;
                1664    :   r_radVal = 363;
                1109    :   r_radVal = 344;
                832     :   r_radVal = 326;
                665     :   r_radVal = 308;
                554     :   r_radVal = 291;
                475     :   r_radVal = 276;
                416     :   r_radVal = 261;
                369     :   r_radVal = 247;
                332     :   r_radVal = 234;
                302     :   r_radVal = 222;
                277     :   r_radVal = 211;
                256     :   r_radVal = 201;
                237     :   r_radVal = 191;
                221     :   r_radVal = 182;
                0       :   r_radVal = 0;
                3584    :   r_radVal = 384;
                1792    :   r_radVal = 366;
                1194    :   r_radVal = 348;
                896     :   r_radVal = 331;
                716     :   r_radVal = 314;
                597     :   r_radVal = 298;
                512     :   r_radVal = 283;
                448     :   r_radVal = 269;
                398     :   r_radVal = 256;
                358     :   r_radVal = 243;
                325     :   r_radVal = 231;
                298     :   r_radVal = 220;
                275     :   r_radVal = 210;
                256     :   r_radVal = 201;
                0       :   r_radVal = 0;
                3840    :   r_radVal = 385;
                1920    :   r_radVal = 368;
                1280    :   r_radVal = 352;
                960     :   r_radVal = 335;
                768     :   r_radVal = 320;
                640     :   r_radVal = 305;
                548     :   r_radVal = 290;
                480     :   r_radVal = 277;
                426     :   r_radVal = 264;
                384     :   r_radVal = 252;
                349     :   r_radVal = 240;
                320     :   r_radVal = 229;
                295     :   r_radVal = 219;
                0       :   r_radVal = 0;
                4096    :   r_radVal = 386;
                2048    :   r_radVal = 370;
                1365    :   r_radVal = 355;
                1024    :   r_radVal = 339;
                819     :   r_radVal = 325;
                682     :   r_radVal = 310;
                585     :   r_radVal = 297;
                512     :   r_radVal = 283;
                455     :   r_radVal = 271;
                409     :   r_radVal = 259;
                372     :   r_radVal = 248;
                0       :   r_radVal = 0;
                4352    :   r_radVal = 387;
                2176    :   r_radVal = 372;
                1450    :   r_radVal = 357;
                1088    :   r_radVal = 343;
                870     :   r_radVal = 329;
                725     :   r_radVal = 315;
                621     :   r_radVal = 302;
                544     :   r_radVal = 290;
                483     :   r_radVal = 277;
                435     :   r_radVal = 266;
                0       :   r_radVal = 0;
                4608    :   r_radVal = 388;
                2304    :   r_radVal = 374;
                1536    :   r_radVal = 360;
                1152    :   r_radVal = 346;
                921     :   r_radVal = 333;
                768     :   r_radVal = 320;
                658     :   r_radVal = 307;
                576     :   r_radVal = 295;
                0       :   r_radVal = 0;
                4864    :   r_radVal = 389;
                2432    :   r_radVal = 375;
                1621    :   r_radVal = 362;
                1216    :   r_radVal = 349;
                972     :   r_radVal = 336;
                810     :   r_radVal = 324;
                default :   r_radVal = r_radVal;
            endcase
        end
    end

    assign o_radVal_q8_8 = r_radVal;
    
endmodule
